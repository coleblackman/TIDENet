VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO conv1_wm_sram_16_100_sky130A
   CLASS BLOCK ;
   SIZE 336.32 BY 356.55 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  114.24 0.0 114.98 1.93 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  127.33 0.0 128.07 1.93 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  140.42 0.0 141.16 1.93 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  154.7 0.0 155.44 1.93 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  167.79 0.0 168.53 1.93 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  180.88 0.0 181.62 1.93 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  192.78 0.0 193.52 1.93 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  207.06 0.0 207.8 1.93 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  220.15 0.0 220.89 1.93 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  233.24 0.0 233.98 1.93 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  246.33 0.0 247.07 1.93 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  259.42 0.0 260.16 1.93 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  272.51 0.0 273.25 1.93 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  285.6 0.0 286.34 1.93 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  298.69 0.0 299.43 1.93 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  311.78 0.0 312.52 1.93 ;
      END
   END din0[15]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  101.15 0.0 101.89 1.93 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 160.65 1.93 161.39 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 161.84 1.93 162.58 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 167.79 1.93 168.53 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 171.36 1.93 172.1 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 176.12 1.93 176.86 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 178.5 1.93 179.24 ;
      END
   END addr0[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 28.56 1.93 29.3 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 32.13 1.93 32.87 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  48.79 0.0 49.53 1.93 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  151.13 0.0 151.87 1.93 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  158.27 0.0 159.01 1.93 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  165.41 0.0 166.15 1.93 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  173.74 0.0 174.48 1.93 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  182.07 0.0 182.81 1.93 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  186.83 0.0 187.57 1.93 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  197.54 0.0 198.28 1.93 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  205.87 0.0 206.61 1.93 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  210.63 0.0 211.37 1.93 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  221.34 0.0 222.08 1.93 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  230.86 0.0 231.6 1.93 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  238.0 0.0 238.74 1.93 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  247.52 0.0 248.26 1.93 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  253.47 0.0 254.21 1.93 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  261.8 0.0 262.54 1.93 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  270.13 0.0 270.87 1.93 ;
      END
   END dout0[15]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  8.33 347.48 330.37 350.6 ;
         LAYER m4 ;
         RECT  8.33 8.33 11.45 350.6 ;
         LAYER m4 ;
         RECT  327.25 8.33 330.37 350.6 ;
         LAYER m3 ;
         RECT  8.33 8.33 330.37 11.45 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m4 ;
         RECT  333.2 2.38 336.32 356.55 ;
         LAYER m3 ;
         RECT  2.38 2.38 336.32 5.5 ;
         LAYER m3 ;
         RECT  2.38 353.43 336.32 356.55 ;
         LAYER m4 ;
         RECT  2.38 2.38 5.5 356.55 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  0.91 0.91 335.41 355.64 ;
   LAYER  m2 ;
      RECT  0.91 0.91 335.41 355.64 ;
   LAYER  m3 ;
      RECT  2.83 159.75 335.41 162.29 ;
      RECT  0.91 163.48 2.83 166.89 ;
      RECT  0.91 169.43 2.83 170.46 ;
      RECT  0.91 173.0 2.83 175.22 ;
      RECT  0.91 30.2 2.83 31.23 ;
      RECT  0.91 33.77 2.83 159.75 ;
      RECT  2.83 162.29 7.43 346.58 ;
      RECT  2.83 346.58 7.43 351.5 ;
      RECT  7.43 162.29 331.27 346.58 ;
      RECT  331.27 162.29 335.41 346.58 ;
      RECT  331.27 346.58 335.41 351.5 ;
      RECT  2.83 7.43 7.43 12.35 ;
      RECT  2.83 12.35 7.43 159.75 ;
      RECT  7.43 12.35 331.27 159.75 ;
      RECT  331.27 7.43 335.41 12.35 ;
      RECT  331.27 12.35 335.41 159.75 ;
      RECT  0.91 0.91 1.48 1.48 ;
      RECT  0.91 1.48 1.48 6.4 ;
      RECT  0.91 6.4 1.48 27.66 ;
      RECT  1.48 0.91 2.83 1.48 ;
      RECT  1.48 6.4 2.83 27.66 ;
      RECT  2.83 0.91 7.43 1.48 ;
      RECT  2.83 6.4 7.43 7.43 ;
      RECT  7.43 0.91 331.27 1.48 ;
      RECT  7.43 6.4 331.27 7.43 ;
      RECT  331.27 0.91 335.41 1.48 ;
      RECT  331.27 6.4 335.41 7.43 ;
      RECT  0.91 180.14 1.48 352.53 ;
      RECT  0.91 352.53 1.48 355.64 ;
      RECT  1.48 180.14 2.83 352.53 ;
      RECT  2.83 351.5 7.43 352.53 ;
      RECT  7.43 351.5 331.27 352.53 ;
      RECT  331.27 351.5 335.41 352.53 ;
   LAYER  m4 ;
      RECT  113.64 2.53 115.58 355.64 ;
      RECT  115.58 0.91 126.73 2.53 ;
      RECT  128.67 0.91 139.82 2.53 ;
      RECT  273.85 0.91 285.0 2.53 ;
      RECT  286.94 0.91 298.09 2.53 ;
      RECT  300.03 0.91 311.18 2.53 ;
      RECT  102.49 0.91 113.64 2.53 ;
      RECT  50.13 0.91 100.55 2.53 ;
      RECT  141.76 0.91 150.53 2.53 ;
      RECT  152.47 0.91 154.1 2.53 ;
      RECT  156.04 0.91 157.67 2.53 ;
      RECT  159.61 0.91 164.81 2.53 ;
      RECT  166.75 0.91 167.19 2.53 ;
      RECT  169.13 0.91 173.14 2.53 ;
      RECT  175.08 0.91 180.28 2.53 ;
      RECT  183.41 0.91 186.23 2.53 ;
      RECT  188.17 0.91 192.18 2.53 ;
      RECT  194.12 0.91 196.94 2.53 ;
      RECT  198.88 0.91 205.27 2.53 ;
      RECT  208.4 0.91 210.03 2.53 ;
      RECT  211.97 0.91 219.55 2.53 ;
      RECT  222.68 0.91 230.26 2.53 ;
      RECT  232.2 0.91 232.64 2.53 ;
      RECT  234.58 0.91 237.4 2.53 ;
      RECT  239.34 0.91 245.73 2.53 ;
      RECT  248.86 0.91 252.87 2.53 ;
      RECT  254.81 0.91 258.82 2.53 ;
      RECT  260.76 0.91 261.2 2.53 ;
      RECT  263.14 0.91 269.53 2.53 ;
      RECT  271.47 0.91 271.91 2.53 ;
      RECT  7.73 2.53 12.05 7.73 ;
      RECT  7.73 351.2 12.05 355.64 ;
      RECT  12.05 2.53 113.64 7.73 ;
      RECT  12.05 7.73 113.64 351.2 ;
      RECT  12.05 351.2 113.64 355.64 ;
      RECT  115.58 2.53 326.65 7.73 ;
      RECT  115.58 7.73 326.65 351.2 ;
      RECT  115.58 351.2 326.65 355.64 ;
      RECT  326.65 2.53 330.97 7.73 ;
      RECT  326.65 351.2 330.97 355.64 ;
      RECT  313.12 0.91 332.6 1.78 ;
      RECT  313.12 1.78 332.6 2.53 ;
      RECT  332.6 0.91 335.41 1.78 ;
      RECT  330.97 2.53 332.6 7.73 ;
      RECT  330.97 7.73 332.6 351.2 ;
      RECT  330.97 351.2 332.6 355.64 ;
      RECT  0.91 0.91 1.78 1.78 ;
      RECT  0.91 1.78 1.78 2.53 ;
      RECT  1.78 0.91 6.1 1.78 ;
      RECT  6.1 0.91 48.19 1.78 ;
      RECT  6.1 1.78 48.19 2.53 ;
      RECT  0.91 2.53 1.78 7.73 ;
      RECT  6.1 2.53 7.73 7.73 ;
      RECT  0.91 7.73 1.78 351.2 ;
      RECT  6.1 7.73 7.73 351.2 ;
      RECT  0.91 351.2 1.78 355.64 ;
      RECT  6.1 351.2 7.73 355.64 ;
   END
END    conv1_wm_sram_16_100_sky130A
END    LIBRARY
