module pool2_layer(
    clk,
    rst,
    blob_din_rdy,
    blob_din_en,
    blob_dout_en,
    blob_dout_rdy,
    blob_dout_eop,
    blob_dout,
    blob_din_eop,
    blob_din);

input clk;
input rst;
output	blob_din_rdy;
input	blob_din_en;
output	blob_dout_en;
input	blob_dout_rdy;
output	blob_dout_eop;
output[11903:0]	blob_dout;
input	blob_din_eop;
input[11903:0]	blob_din;


wire[15:0]	op_dout_72_5;
wire[15:0]	op_dout_72_4;
wire[15:0]	op_dout_72_7;
wire[15:0]	op_dout_72_6;
wire[15:0]	op_dout_72_1;
wire[15:0]	op_dout_72_0;
wire[15:0]	op_dout_72_3;
wire[15:0]	op_dout_72_2;
wire[11903:0]	blob_dout_fifo;
wire[15:0]	op_dout_22_2;
wire[15:0]	op_dout_22_3;
wire[15:0]	op_dout_22_0;
wire[15:0]	op_dout_22_1;
wire[15:0]	op_dout_22_6;
wire[15:0]	op_dout_22_7;
wire[15:0]	op_dout_22_4;
wire[15:0]	op_dout_22_5;
wire[15:0]	op_dout_70_3;
wire[15:0]	op_dout_70_2;
wire[15:0]	op_dout_70_1;
wire[15:0]	op_dout_70_0;
wire[15:0]	op_dout_70_7;
wire[15:0]	op_dout_70_6;
wire[15:0]	op_dout_70_5;
wire[15:0]	op_dout_70_4;
wire[127:0]	op_data_74;
wire[127:0]	op_data_75;
wire[127:0]	op_data_76;
wire[127:0]	op_data_77;
wire[127:0]	op_data_70;
wire[127:0]	op_data_71;
wire[127:0]	op_data_72;
wire[127:0]	op_data_73;
wire[127:0]	op_data_78;
wire[127:0]	op_data_79;
wire[15:0]	op_dout_84_3;
wire[15:0]	op_dout_41_3;
wire[15:0]	op_dout_41_1;
wire[15:0]	op_dout_41_0;
wire[15:0]	op_dout_58_0;
wire[15:0]	op_dout_76_1;
wire[15:0]	op_dout_76_0;
wire[15:0]	op_dout_76_3;
wire[15:0]	op_dout_76_2;
wire[15:0]	op_dout_76_5;
wire[15:0]	op_dout_76_4;
wire[15:0]	op_dout_76_7;
wire[15:0]	op_dout_76_6;
wire[15:0]	op_dout_74_7;
wire[15:0]	op_dout_74_6;
wire[15:0]	op_dout_74_5;
wire[15:0]	op_dout_74_4;
wire[15:0]	op_dout_74_3;
wire[15:0]	op_dout_74_2;
wire[15:0]	op_dout_74_1;
wire[15:0]	op_dout_74_0;
wire[127:0]	op_data_4;
wire[127:0]	op_data_5;
wire[15:0]	op_dout_18_7;
wire[127:0]	op_data_7;
wire[15:0]	op_dout_18_1;
wire[127:0]	op_data_1;
wire[15:0]	op_dout_18_3;
wire[15:0]	op_dout_18_2;
wire[127:0]	op_data_8;
wire[127:0]	op_data_9;
wire[15:0]	op_dout_78_3;
wire[15:0]	op_dout_78_2;
wire[15:0]	op_dout_78_1;
wire[15:0]	op_dout_78_0;
wire[15:0]	op_dout_78_7;
wire[15:0]	op_dout_78_6;
wire[15:0]	op_dout_78_5;
wire[15:0]	op_dout_78_4;
wire[15:0]	op_dout_14_1;
wire[15:0]	op_dout_14_0;
wire[15:0]	op_dout_14_3;
wire[15:0]	op_dout_14_2;
wire[15:0]	op_dout_14_5;
wire[15:0]	op_dout_14_4;
wire[15:0]	op_dout_14_7;
wire[15:0]	op_dout_14_6;
wire[15:0]	op_dout_16_7;
wire[15:0]	op_dout_16_6;
wire[15:0]	op_dout_16_5;
wire[15:0]	op_dout_16_4;
wire[15:0]	op_dout_16_3;
wire[15:0]	op_dout_16_2;
wire[15:0]	op_dout_16_1;
wire[15:0]	op_dout_16_0;
wire[15:0]	op_dout_87_1;
wire[15:0]	op_dout_87_0;
wire[15:0]	op_dout_87_3;
wire[15:0]	op_dout_87_2;
wire[15:0]	op_dout_87_5;
wire[15:0]	op_dout_87_4;
wire[15:0]	op_dout_87_7;
wire[15:0]	op_dout_87_6;
wire[15:0]	op_dout_39_2;
wire[15:0]	op_dout_67_6;
wire[15:0]	op_dout_85_6;
wire[15:0]	op_dout_85_5;
wire[15:0]	op_dout_85_4;
wire[15:0]	op_dout_85_3;
wire[15:0]	op_dout_85_2;
wire[15:0]	op_dout_85_1;
wire[15:0]	op_dout_85_0;
wire[15:0]	op_dout_83_5;
wire[15:0]	op_dout_83_4;
wire[15:0]	op_dout_83_7;
wire[15:0]	op_dout_83_6;
wire[15:0]	op_dout_83_1;
wire[15:0]	op_dout_83_0;
wire[15:0]	op_dout_64_7;
wire[15:0]	op_dout_83_2;
wire[15:0]	op_dout_81_3;
wire[15:0]	op_dout_81_2;
wire[15:0]	op_dout_81_1;
wire[15:0]	op_dout_81_0;
wire[15:0]	op_dout_81_7;
wire[15:0]	op_dout_81_6;
wire[15:0]	op_dout_81_5;
wire[15:0]	op_dout_81_4;
wire[15:0]	op_dout_10_5;
wire[15:0]	op_dout_10_4;
wire[15:0]	op_dout_10_7;
wire[15:0]	op_dout_10_6;
wire[15:0]	op_dout_10_1;
wire[15:0]	op_dout_10_0;
wire[15:0]	op_dout_10_3;
wire[15:0]	op_dout_10_2;
wire[15:0]	op_dout_25_1;
wire[15:0]	op_dout_25_0;
wire[15:0]	op_dout_25_3;
wire[15:0]	op_dout_25_2;
wire[15:0]	op_dout_25_5;
wire[127:0]	op_data_35;
wire[127:0]	op_data_36;
wire[15:0]	op_dout_25_6;
wire[127:0]	op_data_38;
wire[127:0]	op_data_39;
wire[15:0]	op_dout_27_7;
wire[15:0]	op_dout_12_2;
wire[15:0]	op_dout_27_5;
wire[15:0]	op_dout_27_4;
wire[15:0]	op_dout_27_3;
wire[15:0]	op_dout_27_2;
wire[15:0]	op_dout_27_1;
wire[15:0]	op_dout_27_0;
wire[15:0]	op_dout_21_5;
wire[15:0]	op_dout_21_4;
wire[15:0]	op_dout_21_7;
wire[15:0]	op_dout_21_6;
wire[15:0]	op_dout_21_1;
wire[15:0]	op_dout_21_0;
wire[15:0]	op_dout_21_3;
wire[15:0]	op_dout_21_2;
wire[15:0]	op_dout_58_5;
wire[15:0]	op_dout_77_3;
wire[15:0]	op_dout_23_3;
wire[15:0]	op_dout_23_2;
wire[15:0]	op_dout_23_1;
wire[15:0]	op_dout_23_0;
wire[15:0]	op_dout_23_7;
wire[15:0]	op_dout_23_6;
wire[15:0]	op_dout_23_5;
wire[15:0]	op_dout_23_4;
wire[15:0]	op_dout_59_2;
wire	rm_wr_en;
wire[15:0]	op_dout_29_5;
wire[15:0]	op_dout_29_4;
wire[15:0]	op_dout_29_7;
wire[15:0]	op_dout_29_6;
wire[15:0]	op_dout_29_1;
wire[15:0]	op_dout_29_0;
wire[15:0]	op_dout_29_3;
wire[15:0]	op_dout_29_2;
wire[15:0]	op_dout_88_3;
wire[15:0]	op_dout_75_5;
wire[15:0]	op_dout_80_2;
wire[15:0]	op_dout_80_3;
wire[15:0]	op_dout_80_0;
wire[15:0]	op_dout_80_1;
wire[15:0]	op_dout_80_6;
wire[15:0]	op_dout_80_7;
wire[15:0]	op_dout_80_4;
wire[15:0]	op_dout_80_5;
wire[15:0]	op_dout_90_5;
wire[15:0]	op_dout_47_5;
wire[15:0]	op_dout_47_4;
wire[15:0]	op_dout_47_7;
wire[15:0]	op_dout_47_6;
wire[15:0]	op_dout_47_1;
wire[15:0]	op_dout_47_0;
wire[15:0]	op_dout_47_3;
wire[15:0]	op_dout_47_2;
wire[15:0]	op_dout_86_0;
wire[15:0]	op_dout_86_1;
wire[15:0]	op_dout_86_2;
wire[15:0]	op_dout_86_3;
wire[15:0]	op_dout_86_4;
wire[15:0]	op_dout_86_5;
wire[15:0]	op_dout_86_6;
wire[15:0]	op_dout_86_7;
wire[127:0]	op_data_69;
wire[127:0]	op_data_68;
wire[15:0]	op_dout_90_4;
wire[127:0]	op_data_63;
wire[127:0]	op_data_62;
wire[127:0]	op_data_61;
wire[127:0]	op_data_60;
wire[127:0]	op_data_67;
wire[127:0]	op_data_66;
wire[127:0]	op_data_65;
wire[127:0]	op_data_64;
wire[15:0]	op_dout_82_4;
wire[15:0]	op_dout_82_5;
wire[15:0]	op_dout_82_6;
wire[15:0]	op_dout_82_7;
wire[15:0]	op_dout_82_0;
wire[15:0]	op_dout_82_1;
wire[15:0]	op_dout_82_2;
wire[15:0]	op_dout_82_3;
wire[4:0]	rm_rd_addr;
wire[15:0]	op_dout_49_7;
wire[15:0]	op_dout_49_6;
wire[15:0]	op_dout_49_5;
wire[15:0]	op_dout_49_4;
wire[15:0]	op_dout_49_3;
wire[15:0]	op_dout_49_2;
wire[15:0]	op_dout_49_1;
wire[15:0]	op_dout_49_0;
wire[15:0]	op_dout_89_3;
wire[15:0]	op_dout_89_2;
wire[15:0]	op_dout_89_1;
wire[15:0]	op_dout_89_0;
wire[15:0]	op_dout_89_7;
wire[15:0]	op_dout_89_6;
wire[15:0]	op_dout_89_5;
wire[15:0]	op_dout_89_4;
wire[15:0]	op_dout_85_7;
wire[15:0]	op_dout_90_6;
wire[15:0]	op_dout_43_1;
wire[15:0]	op_dout_43_0;
wire[15:0]	op_dout_43_3;
wire[15:0]	op_dout_43_2;
wire[15:0]	op_dout_43_5;
wire[15:0]	op_dout_43_4;
wire[15:0]	op_dout_43_7;
wire[15:0]	op_dout_43_6;
wire[15:0]	op_dout_90_1;
wire[15:0]	op_dout_41_7;
wire[15:0]	op_dout_41_6;
wire[15:0]	op_dout_41_5;
wire[15:0]	op_dout_41_4;
wire[127:0]	op_data_92;
wire[15:0]	op_dout_41_2;
wire[127:0]	op_data_90;
wire[127:0]	op_data_91;
wire[15:0]	op_dout_90_0;
wire[15:0]	op_dout_45_5;
wire[15:0]	op_dout_69_4;
wire[15:0]	op_dout_61_1;
wire[15:0]	op_dout_61_0;
wire[15:0]	op_dout_61_3;
wire[15:0]	op_dout_61_2;
wire[15:0]	op_dout_61_5;
wire[15:0]	op_dout_61_4;
wire[15:0]	op_dout_61_7;
wire[15:0]	op_dout_61_6;
wire[15:0]	op_dout_63_7;
wire[15:0]	op_dout_63_6;
wire[15:0]	op_dout_63_5;
wire[15:0]	op_dout_63_4;
wire[15:0]	op_dout_63_3;
wire[15:0]	op_dout_63_2;
wire[15:0]	op_dout_63_1;
wire[15:0]	op_dout_63_0;
wire[15:0]	op_dout_18_5;
wire[15:0]	op_dout_18_4;
wire[15:0]	op_dout_90_2;
wire[127:0]	op_data_6;
wire[15:0]	op_dout_18_6;
wire[127:0]	op_data_0;
wire[15:0]	op_dout_18_0;
wire[15:0]	op_dout_69_1;
wire[15:0]	op_dout_69_0;
wire[15:0]	op_dout_69_3;
wire[15:0]	op_dout_69_2;
wire[15:0]	op_dout_69_5;
wire[127:0]	op_data_2;
wire[15:0]	op_dout_69_7;
wire[15:0]	op_dout_69_6;
wire[127:0]	op_data_3;
wire[15:0]	op_dout_37_0;
wire[15:0]	op_dout_65_5;
wire[15:0]	op_dout_65_4;
wire[15:0]	op_dout_65_7;
wire[15:0]	op_dout_65_6;
wire[15:0]	op_dout_65_1;
wire[15:0]	op_dout_65_0;
wire[15:0]	op_dout_65_3;
wire[15:0]	op_dout_65_2;
wire[127:0]	op_data_27;
wire[127:0]	op_data_26;
wire[127:0]	op_data_25;
wire[127:0]	op_data_24;
wire[127:0]	op_data_23;
wire[127:0]	op_data_22;
wire[127:0]	op_data_21;
wire[127:0]	op_data_20;
wire[127:0]	op_data_29;
wire[127:0]	op_data_28;
wire[15:0]	op_dout_30_7;
wire[15:0]	op_dout_30_6;
wire[15:0]	op_dout_30_5;
wire[15:0]	op_dout_30_4;
wire[15:0]	op_dout_30_3;
wire[15:0]	op_dout_30_2;
wire[15:0]	op_dout_30_1;
wire[15:0]	op_dout_30_0;
wire[15:0]	op_dout_36_5;
wire[15:0]	op_dout_36_4;
wire[15:0]	op_dout_36_7;
wire[15:0]	op_dout_36_6;
wire[15:0]	op_dout_36_1;
wire[15:0]	op_dout_36_0;
wire[15:0]	op_dout_36_3;
wire[15:0]	op_dout_36_2;
wire[15:0]	op_dout_55_3;
wire	op_din_eop;
wire[15:0]	op_dout_84_6;
wire[4:0]	rm_wr_addr;
wire[127:0]	op_data_52;
wire[127:0]	op_data_53;
wire[127:0]	op_data_50;
wire[127:0]	op_data_51;
wire[127:0]	op_data_56;
wire[127:0]	op_data_57;
wire[127:0]	op_data_54;
wire[127:0]	op_data_55;
wire[127:0]	op_data_58;
wire[127:0]	op_data_59;
wire	op_din_en;
wire[15:0]	op_dout_67_2;
wire[15:0]	op_dout_34_3;
wire[15:0]	op_dout_34_2;
wire[15:0]	op_dout_34_1;
wire[15:0]	op_dout_34_0;
wire[15:0]	op_dout_34_7;
wire[15:0]	op_dout_34_6;
wire[15:0]	op_dout_34_5;
wire[15:0]	op_dout_34_4;
wire[15:0]	op_dout_44_2;
wire[15:0]	op_dout_32_1;
wire[15:0]	op_dout_44_0;
wire[15:0]	op_dout_44_1;
wire[15:0]	op_dout_44_6;
wire[15:0]	op_dout_44_7;
wire[15:0]	op_dout_44_4;
wire[15:0]	op_dout_32_0;
wire[15:0]	op_dout_38_7;
wire[15:0]	op_dout_38_6;
wire[15:0]	op_dout_38_5;
wire[15:0]	op_dout_38_4;
wire[15:0]	op_dout_38_3;
wire[15:0]	op_dout_32_3;
wire[15:0]	op_dout_38_1;
wire[15:0]	op_dout_38_0;
wire[15:0]	op_dout_91_4;
wire[15:0]	op_dout_32_2;
wire[15:0]	op_dout_91_5;
wire[15:0]	op_dout_32_5;
wire[15:0]	op_dout_91_6;
wire[15:0]	op_dout_32_4;
wire[15:0]	op_dout_91_7;
wire[15:0]	op_dout_32_7;
wire[15:0]	op_dout_91_0;
wire[15:0]	op_dout_32_6;
wire[15:0]	op_dout_91_1;
wire[15:0]	op_dout_91_2;
wire[15:0]	op_dout_91_3;
wire[15:0]	op_dout_13_4;
wire[15:0]	op_dout_42_0;
wire[15:0]	op_dout_42_1;
wire[15:0]	op_dout_42_2;
wire[15:0]	op_dout_42_3;
wire[15:0]	op_dout_42_4;
wire[15:0]	op_dout_42_5;
wire[15:0]	op_dout_42_6;
wire[15:0]	op_dout_42_7;
wire[15:0]	op_dout_55_5;
wire[15:0]	op_dout_40_6;
wire[15:0]	op_dout_40_7;
wire[15:0]	op_dout_40_4;
wire[15:0]	op_dout_40_5;
wire[15:0]	op_dout_40_2;
wire[15:0]	op_dout_40_3;
wire[15:0]	op_dout_40_0;
wire[15:0]	op_dout_40_1;
wire[15:0]	op_dout_48_6;
wire[15:0]	op_dout_48_7;
wire[15:0]	op_dout_48_4;
wire[15:0]	op_dout_48_5;
wire[15:0]	op_dout_48_2;
wire[15:0]	op_dout_48_3;
wire[15:0]	op_dout_48_0;
wire[15:0]	op_dout_48_1;
wire[15:0]	op_dout_6_1;
wire[15:0]	op_dout_6_0;
wire[15:0]	op_dout_6_3;
wire[15:0]	op_dout_6_2;
wire[15:0]	op_dout_6_5;
wire[15:0]	op_dout_6_4;
wire[15:0]	op_dout_6_7;
wire[15:0]	op_dout_6_6;
wire[15:0]	op_dout_67_0;
wire[15:0]	op_dout_0_3;
wire[15:0]	op_dout_0_2;
wire[15:0]	op_dout_0_1;
wire[15:0]	op_dout_0_0;
wire[15:0]	op_dout_0_7;
wire[15:0]	op_dout_0_6;
wire[15:0]	op_dout_0_5;
wire[15:0]	op_dout_0_4;
wire[15:0]	op_dout_67_5;
wire[15:0]	op_dout_67_4;
wire[15:0]	op_dout_60_0;
wire[15:0]	op_dout_60_1;
wire[15:0]	op_dout_60_2;
wire[15:0]	op_dout_60_3;
wire[15:0]	op_dout_60_4;
wire[15:0]	op_dout_60_5;
wire[15:0]	op_dout_60_6;
wire[15:0]	op_dout_60_7;
wire[15:0]	op_dout_66_3;
wire[127:0]	op_data_18;
wire[127:0]	op_data_19;
wire[127:0]	op_data_16;
wire[127:0]	op_data_17;
wire[127:0]	op_data_14;
wire[127:0]	op_data_15;
wire[127:0]	op_data_12;
wire[127:0]	op_data_13;
wire[127:0]	op_data_10;
wire[127:0]	op_data_11;
wire[15:0]	op_dout_68_0;
wire[15:0]	op_dout_68_1;
wire[15:0]	op_dout_68_2;
wire[15:0]	op_dout_68_3;
wire[15:0]	op_dout_68_4;
wire[15:0]	op_dout_68_5;
wire[15:0]	op_dout_68_6;
wire[15:0]	op_dout_68_7;
wire[15:0]	op_dout_4_7;
wire[15:0]	op_dout_4_6;
wire[15:0]	op_dout_4_5;
wire[15:0]	op_dout_4_4;
wire[15:0]	op_dout_4_3;
wire[15:0]	op_dout_4_2;
wire[15:0]	op_dout_4_1;
wire[15:0]	op_dout_4_0;
wire[15:0]	op_dout_62_6;
wire[15:0]	op_dout_62_7;
wire[15:0]	op_dout_62_4;
wire[15:0]	op_dout_62_5;
wire[15:0]	op_dout_62_2;
wire[15:0]	op_dout_62_3;
wire[15:0]	op_dout_62_0;
wire[15:0]	op_dout_62_1;
wire[15:0]	op_dout_90_7;
wire[15:0]	op_dout_64_4;
wire[15:0]	op_dout_64_5;
wire[15:0]	op_dout_64_6;
wire[15:0]	op_dout_57_1;
wire[15:0]	op_dout_64_0;
wire[15:0]	op_dout_64_1;
wire[15:0]	op_dout_64_2;
wire[15:0]	op_dout_64_3;
wire[15:0]	op_dout_9_2;
wire[15:0]	op_dout_9_3;
wire[15:0]	op_dout_9_0;
wire[15:0]	op_dout_9_1;
wire[15:0]	op_dout_9_6;
wire[15:0]	op_dout_9_7;
wire[15:0]	op_dout_9_4;
wire[15:0]	op_dout_9_5;
wire[15:0]	op_dout_67_3;
wire[15:0]	op_dout_90_3;
wire[15:0]	op_dout_31_6;
wire[15:0]	op_dout_31_7;
wire[15:0]	op_dout_31_4;
wire[15:0]	op_dout_31_5;
wire[15:0]	op_dout_31_2;
wire[15:0]	op_dout_31_3;
wire[15:0]	op_dout_31_0;
wire[15:0]	op_dout_31_1;
wire[127:0]	op_data_85;
wire[127:0]	op_data_84;
wire[127:0]	op_data_87;
wire[127:0]	op_data_86;
wire[127:0]	op_data_81;
wire[127:0]	op_data_80;
wire[127:0]	op_data_83;
wire[127:0]	op_data_82;
wire[15:0]	op_dout_37_4;
wire[15:0]	op_dout_37_5;
wire[15:0]	op_dout_37_6;
wire[15:0]	op_dout_37_7;
wire[127:0]	op_data_89;
wire[127:0]	op_data_88;
wire[15:0]	op_dout_37_2;
wire[15:0]	op_dout_37_3;
wire[15:0]	op_dout_54_5;
wire[15:0]	op_dout_54_4;
wire[15:0]	op_dout_73_5;
wire[15:0]	op_dout_54_7;
wire[15:0]	op_dout_33_0;
wire[15:0]	op_dout_54_6;
wire[15:0]	op_dout_33_1;
wire[15:0]	op_dout_54_1;
wire[15:0]	op_dout_33_2;
wire[15:0]	op_dout_54_0;
wire[15:0]	op_dout_66_2;
wire[15:0]	op_dout_59_0;
wire[15:0]	op_dout_33_3;
wire[15:0]	op_dout_54_3;
wire[15:0]	op_dout_59_1;
wire[15:0]	op_dout_3_4;
wire[15:0]	op_dout_3_5;
wire[15:0]	op_dout_3_6;
wire[15:0]	op_dout_3_7;
wire[15:0]	op_dout_3_0;
wire[15:0]	op_dout_3_1;
wire[15:0]	op_dout_3_2;
wire[15:0]	op_dout_3_3;
wire[15:0]	op_dout_59_3;
wire[15:0]	op_dout_33_6;
wire[15:0]	op_dout_59_4;
wire[15:0]	op_dout_33_7;
wire[15:0]	op_dout_59_5;
wire[15:0]	op_dout_59_6;
wire[15:0]	op_dout_59_7;
wire[15:0]	op_dout_35_2;
wire[15:0]	op_dout_35_3;
wire[15:0]	op_dout_35_0;
wire[15:0]	op_dout_35_1;
wire[15:0]	op_dout_35_6;
wire[15:0]	op_dout_35_7;
wire[15:0]	op_dout_35_4;
wire[15:0]	op_dout_35_5;
wire[15:0]	op_dout_67_7;
wire[15:0]	op_dout_92_0;
wire[15:0]	op_dout_83_3;
wire[15:0]	op_dout_58_3;
wire[15:0]	op_dout_92_6;
wire[15:0]	op_dout_39_6;
wire[15:0]	op_dout_39_7;
wire[15:0]	op_dout_39_4;
wire[15:0]	op_dout_39_5;
wire[15:0]	op_dout_33_4;
wire[15:0]	op_dout_39_3;
wire[15:0]	op_dout_39_0;
wire[15:0]	op_dout_39_1;
wire[15:0]	op_dout_66_0;
wire[15:0]	op_dout_66_1;
wire[15:0]	op_dout_46_4;
wire[15:0]	op_dout_66_6;
wire[15:0]	op_dout_66_7;
wire[15:0]	op_dout_56_3;
wire[15:0]	op_dout_33_5;
wire[15:0]	op_dout_66_4;
wire[15:0]	op_dout_56_2;
wire	blob_dout_en_fifo;
wire[15:0]	op_dout_66_5;
wire[15:0]	op_dout_56_1;
wire[15:0]	op_dout_56_0;
wire[15:0]	op_dout_56_7;
wire[15:0]	op_dout_56_6;
wire[15:0]	op_dout_56_5;
wire[15:0]	op_dout_56_4;
wire[15:0]	op_dout_7_0;
wire[15:0]	op_dout_7_1;
wire[15:0]	op_dout_7_2;
wire[15:0]	op_dout_7_3;
wire[15:0]	op_dout_7_4;
wire[15:0]	op_dout_7_5;
wire[15:0]	op_dout_7_6;
wire[15:0]	op_dout_7_7;
wire[15:0]	op_dout_1_2;
wire[15:0]	op_dout_1_3;
wire[15:0]	op_dout_1_0;
wire[15:0]	op_dout_1_1;
wire[15:0]	op_dout_1_6;
wire[15:0]	op_dout_1_7;
wire[15:0]	op_dout_1_4;
wire[15:0]	op_dout_1_5;
wire[127:0]	op_data_41;
wire[127:0]	op_data_40;
wire[127:0]	op_data_43;
wire[127:0]	op_data_42;
wire[127:0]	op_data_45;
wire[127:0]	op_data_44;
wire[127:0]	op_data_47;
wire[127:0]	op_data_46;
wire[127:0]	op_data_49;
wire[127:0]	op_data_48;
wire[15:0]	op_dout_37_1;
wire[15:0]	op_dout_26_6;
wire[15:0]	op_dout_46_5;
wire[15:0]	op_dout_58_1;
wire[15:0]	op_dout_26_7;
wire[15:0]	op_dout_13_0;
wire[15:0]	op_dout_26_5;
wire	blob_dout_eop_fifo;
wire[15:0]	op_dout_84_7;
wire[15:0]	op_dout_55_4;
wire[15:0]	op_dout_26_2;
wire[15:0]	op_dout_55_6;
wire[15:0]	op_dout_55_7;
wire[15:0]	op_dout_55_0;
wire[15:0]	op_dout_55_1;
wire[15:0]	op_dout_55_2;
wire[15:0]	op_dout_13_7;
wire[15:0]	op_dout_45_3;
wire[15:0]	op_dout_26_0;
wire[15:0]	op_dout_45_2;
wire[15:0]	op_dout_13_5;
wire[15:0]	op_dout_45_1;
wire[15:0]	op_dout_57_2;
wire[15:0]	op_dout_57_3;
wire[15:0]	op_dout_57_0;
wire[15:0]	op_dout_45_0;
wire[15:0]	op_dout_57_6;
wire[15:0]	op_dout_57_7;
wire[15:0]	op_dout_57_4;
wire[15:0]	op_dout_57_5;
wire[15:0]	op_dout_45_7;
wire[15:0]	op_dout_45_6;
wire[15:0]	op_dout_5_6;
wire[15:0]	op_dout_5_7;
wire[15:0]	op_dout_5_4;
wire[15:0]	op_dout_5_5;
wire[15:0]	op_dout_5_2;
wire[15:0]	op_dout_5_3;
wire[15:0]	op_dout_5_0;
wire[15:0]	op_dout_5_1;
wire[15:0]	op_dout_92_3;
wire[15:0]	op_dout_92_2;
wire[15:0]	op_dout_92_1;
wire[15:0]	op_dout_45_4;
wire[15:0]	op_dout_92_7;
wire[15:0]	op_dout_88_0;
wire[15:0]	op_dout_92_5;
wire[15:0]	op_dout_92_4;
wire[15:0]	op_dout_84_5;
wire[15:0]	op_dout_88_1;
wire[15:0]	op_dout_88_6;
wire[15:0]	op_dout_58_2;
wire[15:0]	op_dout_88_7;
wire[15:0]	op_dout_54_2;
wire[15:0]	op_dout_88_4;
wire[15:0]	op_dout_88_5;
wire[15:0]	op_dout_8_3;
wire[15:0]	op_dout_8_2;
wire[15:0]	op_dout_8_1;
wire[15:0]	op_dout_8_0;
wire[15:0]	op_dout_8_7;
wire[15:0]	op_dout_8_6;
wire[15:0]	op_dout_8_5;
wire[15:0]	op_dout_8_4;
wire[15:0]	op_dout_51_0;
wire[15:0]	op_dout_51_1;
wire[15:0]	op_dout_51_2;
wire[15:0]	op_dout_51_3;
wire[15:0]	op_dout_51_4;
wire[127:0]	op_data_32;
wire[15:0]	op_dout_51_6;
wire[15:0]	op_dout_51_7;
wire[15:0]	op_dout_84_4;
wire[127:0]	op_data_33;
wire[15:0]	op_dout_53_6;
wire[127:0]	op_data_34;
wire[15:0]	op_dout_53_4;
wire[15:0]	op_dout_53_5;
wire[15:0]	op_dout_53_2;
wire[15:0]	op_dout_53_3;
wire[15:0]	op_dout_53_0;
wire[15:0]	op_dout_25_4;
wire[15:0]	op_dout_25_7;
wire[15:0]	op_dout_73_4;
wire[15:0]	op_dout_58_4;
wire[15:0]	op_dout_73_6;
wire[127:0]	op_data_37;
wire[15:0]	op_dout_73_0;
wire[15:0]	op_dout_73_1;
wire[15:0]	op_dout_73_2;
wire[15:0]	op_dout_51_5;
wire[15:0]	op_dout_84_0;
wire[15:0]	op_dout_71_2;
wire[15:0]	op_dout_71_3;
wire[15:0]	op_dout_71_0;
wire[15:0]	op_dout_71_1;
wire[15:0]	op_dout_71_6;
wire[15:0]	op_dout_71_7;
wire[15:0]	op_dout_71_4;
wire[15:0]	op_dout_58_7;
wire[15:0]	op_dout_2_5;
wire[15:0]	op_dout_2_4;
wire[15:0]	op_dout_2_7;
wire[15:0]	op_dout_2_6;
wire[15:0]	op_dout_2_1;
wire[15:0]	op_dout_2_0;
wire[15:0]	op_dout_2_3;
wire[15:0]	op_dout_2_2;
wire[15:0]	op_dout_84_1;
wire[15:0]	op_dout_46_6;
wire[15:0]	op_dout_12_3;
wire[15:0]	op_dout_46_7;
wire[15:0]	op_dout_58_6;
wire[15:0]	op_dout_27_6;
wire[15:0]	op_dout_46_0;
wire[15:0]	op_dout_12_1;
wire[15:0]	op_dout_46_1;
wire[15:0]	op_dout_12_0;
wire[15:0]	op_dout_46_2;
wire[15:0]	op_dout_53_7;
wire[15:0]	op_dout_12_7;
wire[15:0]	op_dout_46_3;
wire[15:0]	op_dout_12_6;
wire[15:0]	op_dout_12_5;
wire[15:0]	op_dout_77_0;
wire[15:0]	op_dout_77_1;
wire[15:0]	op_dout_77_2;
wire[15:0]	op_dout_12_4;
wire[15:0]	op_dout_77_4;
wire[15:0]	op_dout_77_5;
wire[15:0]	op_dout_77_6;
wire[15:0]	op_dout_77_7;
wire[15:0]	op_dout_75_6;
wire[15:0]	op_dout_75_7;
wire[15:0]	op_dout_75_4;
wire[15:0]	op_dout_53_1;
wire[15:0]	op_dout_75_2;
wire[15:0]	op_dout_75_3;
wire[15:0]	op_dout_75_0;
wire[15:0]	op_dout_75_1;
wire[15:0]	op_dout_19_4;
wire[15:0]	op_dout_19_5;
wire[15:0]	op_dout_19_6;
wire[15:0]	op_dout_19_7;
wire[15:0]	op_dout_19_0;
wire[15:0]	op_dout_19_1;
wire[15:0]	op_dout_19_2;
wire[15:0]	op_dout_19_3;
wire[15:0]	op_dout_79_2;
wire[15:0]	op_dout_79_3;
wire[15:0]	op_dout_79_0;
wire[15:0]	op_dout_79_1;
wire[15:0]	op_dout_79_6;
wire[15:0]	op_dout_79_7;
wire[15:0]	op_dout_79_4;
wire[15:0]	op_dout_79_5;
wire[15:0]	op_dout_15_0;
wire[15:0]	op_dout_15_1;
wire[15:0]	op_dout_15_2;
wire[15:0]	op_dout_15_3;
wire[15:0]	op_dout_15_4;
wire[15:0]	op_dout_15_5;
wire[15:0]	op_dout_15_6;
wire[15:0]	op_dout_15_7;
wire[15:0]	op_dout_73_7;
wire[15:0]	op_dout_44_3;
wire[15:0]	op_dout_84_2;
wire[15:0]	op_dout_73_3;
wire[15:0]	op_dout_44_5;
wire[15:0]	op_dout_67_1;
wire[15:0]	op_dout_17_6;
wire[15:0]	op_dout_17_7;
wire[15:0]	op_dout_17_4;
wire[15:0]	op_dout_17_5;
wire[15:0]	op_dout_17_2;
wire[15:0]	op_dout_17_3;
wire[15:0]	op_dout_17_0;
wire[15:0]	op_dout_17_1;
wire[15:0]	op_dout_38_2;
wire[15:0]	op_dout_11_4;
wire[15:0]	op_dout_11_5;
wire[15:0]	op_dout_11_6;
wire[15:0]	op_dout_11_7;
wire[15:0]	op_dout_11_0;
wire[15:0]	op_dout_11_1;
wire[15:0]	op_dout_11_2;
wire[15:0]	op_dout_11_3;
wire[15:0]	op_dout_24_0;
wire[15:0]	op_dout_24_1;
wire[15:0]	op_dout_24_2;
wire[15:0]	op_dout_24_3;
wire[15:0]	op_dout_24_4;
wire[15:0]	op_dout_24_5;
wire[15:0]	op_dout_24_6;
wire[15:0]	op_dout_24_7;
wire[15:0]	op_dout_13_2;
wire[15:0]	op_dout_13_3;
wire[15:0]	op_dout_26_4;
wire[15:0]	op_dout_13_1;
wire[15:0]	op_dout_13_6;
wire[15:0]	op_dout_26_3;
wire[127:0]	op_data_30;
wire[15:0]	op_dout_26_1;
wire[15:0]	op_dout_20_4;
wire[15:0]	op_dout_20_5;
wire[15:0]	op_dout_20_6;
wire[15:0]	op_dout_20_7;
wire[15:0]	op_dout_20_0;
wire[15:0]	op_dout_20_1;
wire[15:0]	op_dout_20_2;
wire[15:0]	op_dout_20_3;
wire[15:0]	op_dout_28_4;
wire[15:0]	op_dout_28_5;
wire[15:0]	op_dout_28_6;
wire[15:0]	op_dout_28_7;
wire[15:0]	op_dout_28_0;
wire[15:0]	op_dout_28_1;
wire[15:0]	op_dout_28_2;
wire[15:0]	op_dout_28_3;
wire[127:0]	op_data_31;
wire[15:0]	op_dout_50_1;
wire[15:0]	op_dout_50_0;
wire[15:0]	op_dout_50_3;
wire[15:0]	op_dout_50_2;
wire[15:0]	op_dout_50_5;
wire[15:0]	op_dout_50_4;
wire[15:0]	op_dout_50_7;
wire[15:0]	op_dout_50_6;
wire[15:0]	op_dout_71_5;
wire[15:0]	op_dout_52_7;
wire[15:0]	op_dout_52_6;
wire[15:0]	op_dout_52_5;
wire[15:0]	op_dout_52_4;
wire[15:0]	op_dout_52_3;
wire[15:0]	op_dout_52_2;
wire[15:0]	op_dout_52_1;
wire[15:0]	op_dout_52_0;
wire[15:0]	op_dout_88_2;


controller_v2_a #(
.DB_W_IN (8),
.DB_H_IN (8),
.DB_C_IN (8),
.DB_W_OUT (4),
.DB_H_OUT (4),
.DB_C_OUT (8),
.WB_W (2),
.WB_H (2),
.WB_K (8),
.RM_WR_ADDR_WIDTH (5),
.RM_WR_NUM_PER_CHANNEL (1),
.RM_WR_STRIDE (1),
.RM_RING_LENGTH (4),
.RM_RD_PHY_ADDR_JUMP (2),
.RM_RD_ADDR_WIDTH (5),
.KPF (8),
.STRIDE_H (2),
.STRIDE_W (2),
.PAD (0),
.DATA_ACCESS_DELAY (5),
.OP_DELAY (1))
u_controller(
.clk(clk),
.rst(rst),
.rm_wr_en(rm_wr_en), 
.rm_wr_addr(rm_wr_addr),
.rm_rd_addr(rm_rd_addr),
.op_din_eop(op_din_eop),
.op_din_en(op_din_en),
.blob_din_rdy(blob_din_rdy),
.blob_din_en(blob_din_en), 
.blob_din_eop(blob_din_eop),
.blob_dout_rdy(blob_dout_rdy),
.blob_dout_en(blob_dout_en_fifo),
.blob_dout_eop(blob_dout_eop_fifo));

pool2_rm_ram u_pool2_rm_ram_0(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[127:0]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_0));

pool2_rm_ram u_pool2_rm_ram_1(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[255:128]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_1));

pool2_rm_ram u_pool2_rm_ram_2(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[383:256]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_2));

pool2_rm_ram u_pool2_rm_ram_3(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[511:384]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_3));

pool2_rm_ram u_pool2_rm_ram_4(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[639:512]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_4));

pool2_rm_ram u_pool2_rm_ram_5(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[767:640]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_5));

pool2_rm_ram u_pool2_rm_ram_6(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[895:768]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_6));

pool2_rm_ram u_pool2_rm_ram_7(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[1023:896]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_7));

pool2_rm_ram u_pool2_rm_ram_8(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[1151:1024]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_8));

pool2_rm_ram u_pool2_rm_ram_9(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[1279:1152]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_9));

pool2_rm_ram u_pool2_rm_ram_10(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[1407:1280]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_10));

pool2_rm_ram u_pool2_rm_ram_11(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[1535:1408]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_11));

pool2_rm_ram u_pool2_rm_ram_12(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[1663:1536]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_12));

pool2_rm_ram u_pool2_rm_ram_13(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[1791:1664]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_13));

pool2_rm_ram u_pool2_rm_ram_14(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[1919:1792]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_14));

pool2_rm_ram u_pool2_rm_ram_15(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[2047:1920]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_15));

pool2_rm_ram u_pool2_rm_ram_16(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[2175:2048]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_16));

pool2_rm_ram u_pool2_rm_ram_17(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[2303:2176]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_17));

pool2_rm_ram u_pool2_rm_ram_18(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[2431:2304]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_18));

pool2_rm_ram u_pool2_rm_ram_19(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[2559:2432]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_19));

pool2_rm_ram u_pool2_rm_ram_20(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[2687:2560]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_20));

pool2_rm_ram u_pool2_rm_ram_21(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[2815:2688]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_21));

pool2_rm_ram u_pool2_rm_ram_22(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[2943:2816]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_22));

pool2_rm_ram u_pool2_rm_ram_23(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[3071:2944]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_23));

pool2_rm_ram u_pool2_rm_ram_24(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[3199:3072]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_24));

pool2_rm_ram u_pool2_rm_ram_25(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[3327:3200]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_25));

pool2_rm_ram u_pool2_rm_ram_26(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[3455:3328]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_26));

pool2_rm_ram u_pool2_rm_ram_27(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[3583:3456]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_27));

pool2_rm_ram u_pool2_rm_ram_28(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[3711:3584]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_28));

pool2_rm_ram u_pool2_rm_ram_29(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[3839:3712]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_29));

pool2_rm_ram u_pool2_rm_ram_30(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[3967:3840]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_30));

pool2_rm_ram u_pool2_rm_ram_31(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[4095:3968]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_31));

pool2_rm_ram u_pool2_rm_ram_32(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[4223:4096]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_32));

pool2_rm_ram u_pool2_rm_ram_33(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[4351:4224]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_33));

pool2_rm_ram u_pool2_rm_ram_34(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[4479:4352]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_34));

pool2_rm_ram u_pool2_rm_ram_35(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[4607:4480]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_35));

pool2_rm_ram u_pool2_rm_ram_36(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[4735:4608]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_36));

pool2_rm_ram u_pool2_rm_ram_37(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[4863:4736]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_37));

pool2_rm_ram u_pool2_rm_ram_38(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[4991:4864]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_38));

pool2_rm_ram u_pool2_rm_ram_39(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[5119:4992]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_39));

pool2_rm_ram u_pool2_rm_ram_40(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[5247:5120]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_40));

pool2_rm_ram u_pool2_rm_ram_41(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[5375:5248]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_41));

pool2_rm_ram u_pool2_rm_ram_42(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[5503:5376]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_42));

pool2_rm_ram u_pool2_rm_ram_43(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[5631:5504]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_43));

pool2_rm_ram u_pool2_rm_ram_44(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[5759:5632]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_44));

pool2_rm_ram u_pool2_rm_ram_45(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[5887:5760]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_45));

pool2_rm_ram u_pool2_rm_ram_46(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[6015:5888]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_46));

pool2_rm_ram u_pool2_rm_ram_47(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[6143:6016]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_47));

pool2_rm_ram u_pool2_rm_ram_48(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[6271:6144]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_48));

pool2_rm_ram u_pool2_rm_ram_49(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[6399:6272]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_49));

pool2_rm_ram u_pool2_rm_ram_50(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[6527:6400]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_50));

pool2_rm_ram u_pool2_rm_ram_51(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[6655:6528]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_51));

pool2_rm_ram u_pool2_rm_ram_52(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[6783:6656]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_52));

pool2_rm_ram u_pool2_rm_ram_53(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[6911:6784]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_53));

pool2_rm_ram u_pool2_rm_ram_54(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[7039:6912]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_54));

pool2_rm_ram u_pool2_rm_ram_55(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[7167:7040]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_55));

pool2_rm_ram u_pool2_rm_ram_56(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[7295:7168]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_56));

pool2_rm_ram u_pool2_rm_ram_57(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[7423:7296]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_57));

pool2_rm_ram u_pool2_rm_ram_58(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[7551:7424]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_58));

pool2_rm_ram u_pool2_rm_ram_59(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[7679:7552]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_59));

pool2_rm_ram u_pool2_rm_ram_60(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[7807:7680]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_60));

pool2_rm_ram u_pool2_rm_ram_61(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[7935:7808]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_61));

pool2_rm_ram u_pool2_rm_ram_62(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[8063:7936]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_62));

pool2_rm_ram u_pool2_rm_ram_63(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[8191:8064]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_63));

pool2_rm_ram u_pool2_rm_ram_64(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[8319:8192]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_64));

pool2_rm_ram u_pool2_rm_ram_65(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[8447:8320]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_65));

pool2_rm_ram u_pool2_rm_ram_66(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[8575:8448]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_66));

pool2_rm_ram u_pool2_rm_ram_67(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[8703:8576]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_67));

pool2_rm_ram u_pool2_rm_ram_68(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[8831:8704]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_68));

pool2_rm_ram u_pool2_rm_ram_69(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[8959:8832]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_69));

pool2_rm_ram u_pool2_rm_ram_70(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[9087:8960]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_70));

pool2_rm_ram u_pool2_rm_ram_71(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[9215:9088]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_71));

pool2_rm_ram u_pool2_rm_ram_72(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[9343:9216]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_72));

pool2_rm_ram u_pool2_rm_ram_73(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[9471:9344]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_73));

pool2_rm_ram u_pool2_rm_ram_74(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[9599:9472]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_74));

pool2_rm_ram u_pool2_rm_ram_75(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[9727:9600]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_75));

pool2_rm_ram u_pool2_rm_ram_76(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[9855:9728]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_76));

pool2_rm_ram u_pool2_rm_ram_77(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[9983:9856]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_77));

pool2_rm_ram u_pool2_rm_ram_78(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[10111:9984]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_78));

pool2_rm_ram u_pool2_rm_ram_79(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[10239:10112]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_79));

pool2_rm_ram u_pool2_rm_ram_80(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[10367:10240]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_80));

pool2_rm_ram u_pool2_rm_ram_81(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[10495:10368]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_81));

pool2_rm_ram u_pool2_rm_ram_82(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[10623:10496]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_82));

pool2_rm_ram u_pool2_rm_ram_83(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[10751:10624]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_83));

pool2_rm_ram u_pool2_rm_ram_84(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[10879:10752]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_84));

pool2_rm_ram u_pool2_rm_ram_85(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[11007:10880]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_85));

pool2_rm_ram u_pool2_rm_ram_86(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[11135:11008]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_86));

pool2_rm_ram u_pool2_rm_ram_87(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[11263:11136]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_87));

pool2_rm_ram u_pool2_rm_ram_88(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[11391:11264]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_88));

pool2_rm_ram u_pool2_rm_ram_89(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[11519:11392]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_89));

pool2_rm_ram u_pool2_rm_ram_90(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[11647:11520]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_90));

pool2_rm_ram u_pool2_rm_ram_91(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[11775:11648]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_91));

pool2_rm_ram u_pool2_rm_ram_92(
.clka(clk),
.wea(rm_wr_en),
.addra(rm_wr_addr),
.dina(blob_din[11903:11776]),
.clkb(clk),
.addrb(rm_rd_addr),
.doutb(op_data_92));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_0_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_0[15:0]),
.op_dout(op_dout_0_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_0_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_0[31:16]),
.op_dout(op_dout_0_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_0_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_0[47:32]),
.op_dout(op_dout_0_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_0_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_0[63:48]),
.op_dout(op_dout_0_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_0_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_0[79:64]),
.op_dout(op_dout_0_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_0_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_0[95:80]),
.op_dout(op_dout_0_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_0_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_0[111:96]),
.op_dout(op_dout_0_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_0_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_0[127:112]),
.op_dout(op_dout_0_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_1_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_1[15:0]),
.op_dout(op_dout_1_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_1_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_1[31:16]),
.op_dout(op_dout_1_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_1_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_1[47:32]),
.op_dout(op_dout_1_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_1_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_1[63:48]),
.op_dout(op_dout_1_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_1_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_1[79:64]),
.op_dout(op_dout_1_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_1_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_1[95:80]),
.op_dout(op_dout_1_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_1_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_1[111:96]),
.op_dout(op_dout_1_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_1_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_1[127:112]),
.op_dout(op_dout_1_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_2_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_2[15:0]),
.op_dout(op_dout_2_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_2_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_2[31:16]),
.op_dout(op_dout_2_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_2_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_2[47:32]),
.op_dout(op_dout_2_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_2_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_2[63:48]),
.op_dout(op_dout_2_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_2_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_2[79:64]),
.op_dout(op_dout_2_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_2_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_2[95:80]),
.op_dout(op_dout_2_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_2_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_2[111:96]),
.op_dout(op_dout_2_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_2_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_2[127:112]),
.op_dout(op_dout_2_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_3_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_3[15:0]),
.op_dout(op_dout_3_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_3_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_3[31:16]),
.op_dout(op_dout_3_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_3_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_3[47:32]),
.op_dout(op_dout_3_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_3_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_3[63:48]),
.op_dout(op_dout_3_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_3_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_3[79:64]),
.op_dout(op_dout_3_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_3_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_3[95:80]),
.op_dout(op_dout_3_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_3_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_3[111:96]),
.op_dout(op_dout_3_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_3_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_3[127:112]),
.op_dout(op_dout_3_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_4_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_4[15:0]),
.op_dout(op_dout_4_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_4_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_4[31:16]),
.op_dout(op_dout_4_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_4_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_4[47:32]),
.op_dout(op_dout_4_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_4_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_4[63:48]),
.op_dout(op_dout_4_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_4_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_4[79:64]),
.op_dout(op_dout_4_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_4_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_4[95:80]),
.op_dout(op_dout_4_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_4_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_4[111:96]),
.op_dout(op_dout_4_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_4_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_4[127:112]),
.op_dout(op_dout_4_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_5_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_5[15:0]),
.op_dout(op_dout_5_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_5_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_5[31:16]),
.op_dout(op_dout_5_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_5_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_5[47:32]),
.op_dout(op_dout_5_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_5_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_5[63:48]),
.op_dout(op_dout_5_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_5_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_5[79:64]),
.op_dout(op_dout_5_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_5_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_5[95:80]),
.op_dout(op_dout_5_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_5_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_5[111:96]),
.op_dout(op_dout_5_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_5_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_5[127:112]),
.op_dout(op_dout_5_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_6_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_6[15:0]),
.op_dout(op_dout_6_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_6_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_6[31:16]),
.op_dout(op_dout_6_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_6_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_6[47:32]),
.op_dout(op_dout_6_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_6_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_6[63:48]),
.op_dout(op_dout_6_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_6_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_6[79:64]),
.op_dout(op_dout_6_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_6_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_6[95:80]),
.op_dout(op_dout_6_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_6_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_6[111:96]),
.op_dout(op_dout_6_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_6_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_6[127:112]),
.op_dout(op_dout_6_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_7_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_7[15:0]),
.op_dout(op_dout_7_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_7_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_7[31:16]),
.op_dout(op_dout_7_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_7_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_7[47:32]),
.op_dout(op_dout_7_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_7_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_7[63:48]),
.op_dout(op_dout_7_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_7_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_7[79:64]),
.op_dout(op_dout_7_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_7_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_7[95:80]),
.op_dout(op_dout_7_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_7_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_7[111:96]),
.op_dout(op_dout_7_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_7_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_7[127:112]),
.op_dout(op_dout_7_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_8_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_8[15:0]),
.op_dout(op_dout_8_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_8_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_8[31:16]),
.op_dout(op_dout_8_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_8_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_8[47:32]),
.op_dout(op_dout_8_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_8_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_8[63:48]),
.op_dout(op_dout_8_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_8_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_8[79:64]),
.op_dout(op_dout_8_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_8_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_8[95:80]),
.op_dout(op_dout_8_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_8_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_8[111:96]),
.op_dout(op_dout_8_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_8_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_8[127:112]),
.op_dout(op_dout_8_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_9_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_9[15:0]),
.op_dout(op_dout_9_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_9_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_9[31:16]),
.op_dout(op_dout_9_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_9_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_9[47:32]),
.op_dout(op_dout_9_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_9_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_9[63:48]),
.op_dout(op_dout_9_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_9_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_9[79:64]),
.op_dout(op_dout_9_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_9_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_9[95:80]),
.op_dout(op_dout_9_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_9_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_9[111:96]),
.op_dout(op_dout_9_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_9_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_9[127:112]),
.op_dout(op_dout_9_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_10_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_10[15:0]),
.op_dout(op_dout_10_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_10_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_10[31:16]),
.op_dout(op_dout_10_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_10_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_10[47:32]),
.op_dout(op_dout_10_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_10_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_10[63:48]),
.op_dout(op_dout_10_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_10_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_10[79:64]),
.op_dout(op_dout_10_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_10_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_10[95:80]),
.op_dout(op_dout_10_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_10_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_10[111:96]),
.op_dout(op_dout_10_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_10_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_10[127:112]),
.op_dout(op_dout_10_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_11_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_11[15:0]),
.op_dout(op_dout_11_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_11_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_11[31:16]),
.op_dout(op_dout_11_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_11_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_11[47:32]),
.op_dout(op_dout_11_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_11_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_11[63:48]),
.op_dout(op_dout_11_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_11_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_11[79:64]),
.op_dout(op_dout_11_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_11_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_11[95:80]),
.op_dout(op_dout_11_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_11_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_11[111:96]),
.op_dout(op_dout_11_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_11_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_11[127:112]),
.op_dout(op_dout_11_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_12_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_12[15:0]),
.op_dout(op_dout_12_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_12_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_12[31:16]),
.op_dout(op_dout_12_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_12_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_12[47:32]),
.op_dout(op_dout_12_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_12_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_12[63:48]),
.op_dout(op_dout_12_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_12_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_12[79:64]),
.op_dout(op_dout_12_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_12_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_12[95:80]),
.op_dout(op_dout_12_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_12_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_12[111:96]),
.op_dout(op_dout_12_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_12_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_12[127:112]),
.op_dout(op_dout_12_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_13_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_13[15:0]),
.op_dout(op_dout_13_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_13_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_13[31:16]),
.op_dout(op_dout_13_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_13_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_13[47:32]),
.op_dout(op_dout_13_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_13_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_13[63:48]),
.op_dout(op_dout_13_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_13_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_13[79:64]),
.op_dout(op_dout_13_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_13_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_13[95:80]),
.op_dout(op_dout_13_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_13_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_13[111:96]),
.op_dout(op_dout_13_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_13_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_13[127:112]),
.op_dout(op_dout_13_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_14_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_14[15:0]),
.op_dout(op_dout_14_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_14_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_14[31:16]),
.op_dout(op_dout_14_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_14_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_14[47:32]),
.op_dout(op_dout_14_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_14_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_14[63:48]),
.op_dout(op_dout_14_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_14_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_14[79:64]),
.op_dout(op_dout_14_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_14_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_14[95:80]),
.op_dout(op_dout_14_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_14_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_14[111:96]),
.op_dout(op_dout_14_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_14_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_14[127:112]),
.op_dout(op_dout_14_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_15_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_15[15:0]),
.op_dout(op_dout_15_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_15_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_15[31:16]),
.op_dout(op_dout_15_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_15_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_15[47:32]),
.op_dout(op_dout_15_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_15_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_15[63:48]),
.op_dout(op_dout_15_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_15_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_15[79:64]),
.op_dout(op_dout_15_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_15_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_15[95:80]),
.op_dout(op_dout_15_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_15_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_15[111:96]),
.op_dout(op_dout_15_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_15_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_15[127:112]),
.op_dout(op_dout_15_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_16_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_16[15:0]),
.op_dout(op_dout_16_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_16_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_16[31:16]),
.op_dout(op_dout_16_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_16_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_16[47:32]),
.op_dout(op_dout_16_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_16_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_16[63:48]),
.op_dout(op_dout_16_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_16_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_16[79:64]),
.op_dout(op_dout_16_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_16_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_16[95:80]),
.op_dout(op_dout_16_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_16_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_16[111:96]),
.op_dout(op_dout_16_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_16_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_16[127:112]),
.op_dout(op_dout_16_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_17_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_17[15:0]),
.op_dout(op_dout_17_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_17_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_17[31:16]),
.op_dout(op_dout_17_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_17_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_17[47:32]),
.op_dout(op_dout_17_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_17_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_17[63:48]),
.op_dout(op_dout_17_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_17_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_17[79:64]),
.op_dout(op_dout_17_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_17_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_17[95:80]),
.op_dout(op_dout_17_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_17_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_17[111:96]),
.op_dout(op_dout_17_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_17_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_17[127:112]),
.op_dout(op_dout_17_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_18_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_18[15:0]),
.op_dout(op_dout_18_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_18_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_18[31:16]),
.op_dout(op_dout_18_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_18_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_18[47:32]),
.op_dout(op_dout_18_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_18_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_18[63:48]),
.op_dout(op_dout_18_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_18_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_18[79:64]),
.op_dout(op_dout_18_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_18_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_18[95:80]),
.op_dout(op_dout_18_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_18_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_18[111:96]),
.op_dout(op_dout_18_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_18_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_18[127:112]),
.op_dout(op_dout_18_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_19_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_19[15:0]),
.op_dout(op_dout_19_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_19_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_19[31:16]),
.op_dout(op_dout_19_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_19_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_19[47:32]),
.op_dout(op_dout_19_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_19_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_19[63:48]),
.op_dout(op_dout_19_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_19_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_19[79:64]),
.op_dout(op_dout_19_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_19_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_19[95:80]),
.op_dout(op_dout_19_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_19_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_19[111:96]),
.op_dout(op_dout_19_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_19_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_19[127:112]),
.op_dout(op_dout_19_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_20_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_20[15:0]),
.op_dout(op_dout_20_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_20_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_20[31:16]),
.op_dout(op_dout_20_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_20_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_20[47:32]),
.op_dout(op_dout_20_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_20_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_20[63:48]),
.op_dout(op_dout_20_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_20_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_20[79:64]),
.op_dout(op_dout_20_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_20_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_20[95:80]),
.op_dout(op_dout_20_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_20_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_20[111:96]),
.op_dout(op_dout_20_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_20_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_20[127:112]),
.op_dout(op_dout_20_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_21_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_21[15:0]),
.op_dout(op_dout_21_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_21_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_21[31:16]),
.op_dout(op_dout_21_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_21_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_21[47:32]),
.op_dout(op_dout_21_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_21_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_21[63:48]),
.op_dout(op_dout_21_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_21_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_21[79:64]),
.op_dout(op_dout_21_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_21_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_21[95:80]),
.op_dout(op_dout_21_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_21_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_21[111:96]),
.op_dout(op_dout_21_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_21_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_21[127:112]),
.op_dout(op_dout_21_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_22_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_22[15:0]),
.op_dout(op_dout_22_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_22_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_22[31:16]),
.op_dout(op_dout_22_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_22_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_22[47:32]),
.op_dout(op_dout_22_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_22_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_22[63:48]),
.op_dout(op_dout_22_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_22_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_22[79:64]),
.op_dout(op_dout_22_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_22_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_22[95:80]),
.op_dout(op_dout_22_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_22_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_22[111:96]),
.op_dout(op_dout_22_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_22_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_22[127:112]),
.op_dout(op_dout_22_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_23_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_23[15:0]),
.op_dout(op_dout_23_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_23_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_23[31:16]),
.op_dout(op_dout_23_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_23_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_23[47:32]),
.op_dout(op_dout_23_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_23_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_23[63:48]),
.op_dout(op_dout_23_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_23_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_23[79:64]),
.op_dout(op_dout_23_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_23_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_23[95:80]),
.op_dout(op_dout_23_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_23_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_23[111:96]),
.op_dout(op_dout_23_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_23_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_23[127:112]),
.op_dout(op_dout_23_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_24_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_24[15:0]),
.op_dout(op_dout_24_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_24_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_24[31:16]),
.op_dout(op_dout_24_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_24_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_24[47:32]),
.op_dout(op_dout_24_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_24_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_24[63:48]),
.op_dout(op_dout_24_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_24_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_24[79:64]),
.op_dout(op_dout_24_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_24_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_24[95:80]),
.op_dout(op_dout_24_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_24_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_24[111:96]),
.op_dout(op_dout_24_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_24_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_24[127:112]),
.op_dout(op_dout_24_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_25_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_25[15:0]),
.op_dout(op_dout_25_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_25_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_25[31:16]),
.op_dout(op_dout_25_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_25_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_25[47:32]),
.op_dout(op_dout_25_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_25_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_25[63:48]),
.op_dout(op_dout_25_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_25_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_25[79:64]),
.op_dout(op_dout_25_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_25_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_25[95:80]),
.op_dout(op_dout_25_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_25_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_25[111:96]),
.op_dout(op_dout_25_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_25_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_25[127:112]),
.op_dout(op_dout_25_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_26_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_26[15:0]),
.op_dout(op_dout_26_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_26_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_26[31:16]),
.op_dout(op_dout_26_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_26_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_26[47:32]),
.op_dout(op_dout_26_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_26_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_26[63:48]),
.op_dout(op_dout_26_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_26_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_26[79:64]),
.op_dout(op_dout_26_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_26_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_26[95:80]),
.op_dout(op_dout_26_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_26_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_26[111:96]),
.op_dout(op_dout_26_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_26_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_26[127:112]),
.op_dout(op_dout_26_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_27_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_27[15:0]),
.op_dout(op_dout_27_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_27_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_27[31:16]),
.op_dout(op_dout_27_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_27_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_27[47:32]),
.op_dout(op_dout_27_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_27_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_27[63:48]),
.op_dout(op_dout_27_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_27_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_27[79:64]),
.op_dout(op_dout_27_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_27_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_27[95:80]),
.op_dout(op_dout_27_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_27_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_27[111:96]),
.op_dout(op_dout_27_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_27_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_27[127:112]),
.op_dout(op_dout_27_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_28_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_28[15:0]),
.op_dout(op_dout_28_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_28_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_28[31:16]),
.op_dout(op_dout_28_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_28_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_28[47:32]),
.op_dout(op_dout_28_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_28_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_28[63:48]),
.op_dout(op_dout_28_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_28_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_28[79:64]),
.op_dout(op_dout_28_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_28_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_28[95:80]),
.op_dout(op_dout_28_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_28_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_28[111:96]),
.op_dout(op_dout_28_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_28_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_28[127:112]),
.op_dout(op_dout_28_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_29_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_29[15:0]),
.op_dout(op_dout_29_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_29_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_29[31:16]),
.op_dout(op_dout_29_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_29_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_29[47:32]),
.op_dout(op_dout_29_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_29_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_29[63:48]),
.op_dout(op_dout_29_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_29_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_29[79:64]),
.op_dout(op_dout_29_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_29_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_29[95:80]),
.op_dout(op_dout_29_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_29_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_29[111:96]),
.op_dout(op_dout_29_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_29_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_29[127:112]),
.op_dout(op_dout_29_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_30_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_30[15:0]),
.op_dout(op_dout_30_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_30_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_30[31:16]),
.op_dout(op_dout_30_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_30_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_30[47:32]),
.op_dout(op_dout_30_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_30_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_30[63:48]),
.op_dout(op_dout_30_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_30_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_30[79:64]),
.op_dout(op_dout_30_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_30_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_30[95:80]),
.op_dout(op_dout_30_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_30_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_30[111:96]),
.op_dout(op_dout_30_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_30_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_30[127:112]),
.op_dout(op_dout_30_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_31_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_31[15:0]),
.op_dout(op_dout_31_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_31_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_31[31:16]),
.op_dout(op_dout_31_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_31_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_31[47:32]),
.op_dout(op_dout_31_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_31_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_31[63:48]),
.op_dout(op_dout_31_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_31_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_31[79:64]),
.op_dout(op_dout_31_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_31_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_31[95:80]),
.op_dout(op_dout_31_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_31_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_31[111:96]),
.op_dout(op_dout_31_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_31_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_31[127:112]),
.op_dout(op_dout_31_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_32_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_32[15:0]),
.op_dout(op_dout_32_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_32_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_32[31:16]),
.op_dout(op_dout_32_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_32_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_32[47:32]),
.op_dout(op_dout_32_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_32_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_32[63:48]),
.op_dout(op_dout_32_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_32_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_32[79:64]),
.op_dout(op_dout_32_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_32_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_32[95:80]),
.op_dout(op_dout_32_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_32_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_32[111:96]),
.op_dout(op_dout_32_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_32_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_32[127:112]),
.op_dout(op_dout_32_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_33_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_33[15:0]),
.op_dout(op_dout_33_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_33_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_33[31:16]),
.op_dout(op_dout_33_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_33_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_33[47:32]),
.op_dout(op_dout_33_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_33_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_33[63:48]),
.op_dout(op_dout_33_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_33_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_33[79:64]),
.op_dout(op_dout_33_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_33_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_33[95:80]),
.op_dout(op_dout_33_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_33_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_33[111:96]),
.op_dout(op_dout_33_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_33_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_33[127:112]),
.op_dout(op_dout_33_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_34_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_34[15:0]),
.op_dout(op_dout_34_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_34_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_34[31:16]),
.op_dout(op_dout_34_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_34_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_34[47:32]),
.op_dout(op_dout_34_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_34_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_34[63:48]),
.op_dout(op_dout_34_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_34_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_34[79:64]),
.op_dout(op_dout_34_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_34_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_34[95:80]),
.op_dout(op_dout_34_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_34_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_34[111:96]),
.op_dout(op_dout_34_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_34_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_34[127:112]),
.op_dout(op_dout_34_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_35_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_35[15:0]),
.op_dout(op_dout_35_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_35_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_35[31:16]),
.op_dout(op_dout_35_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_35_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_35[47:32]),
.op_dout(op_dout_35_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_35_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_35[63:48]),
.op_dout(op_dout_35_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_35_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_35[79:64]),
.op_dout(op_dout_35_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_35_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_35[95:80]),
.op_dout(op_dout_35_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_35_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_35[111:96]),
.op_dout(op_dout_35_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_35_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_35[127:112]),
.op_dout(op_dout_35_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_36_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_36[15:0]),
.op_dout(op_dout_36_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_36_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_36[31:16]),
.op_dout(op_dout_36_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_36_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_36[47:32]),
.op_dout(op_dout_36_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_36_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_36[63:48]),
.op_dout(op_dout_36_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_36_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_36[79:64]),
.op_dout(op_dout_36_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_36_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_36[95:80]),
.op_dout(op_dout_36_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_36_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_36[111:96]),
.op_dout(op_dout_36_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_36_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_36[127:112]),
.op_dout(op_dout_36_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_37_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_37[15:0]),
.op_dout(op_dout_37_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_37_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_37[31:16]),
.op_dout(op_dout_37_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_37_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_37[47:32]),
.op_dout(op_dout_37_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_37_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_37[63:48]),
.op_dout(op_dout_37_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_37_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_37[79:64]),
.op_dout(op_dout_37_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_37_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_37[95:80]),
.op_dout(op_dout_37_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_37_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_37[111:96]),
.op_dout(op_dout_37_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_37_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_37[127:112]),
.op_dout(op_dout_37_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_38_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_38[15:0]),
.op_dout(op_dout_38_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_38_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_38[31:16]),
.op_dout(op_dout_38_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_38_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_38[47:32]),
.op_dout(op_dout_38_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_38_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_38[63:48]),
.op_dout(op_dout_38_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_38_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_38[79:64]),
.op_dout(op_dout_38_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_38_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_38[95:80]),
.op_dout(op_dout_38_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_38_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_38[111:96]),
.op_dout(op_dout_38_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_38_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_38[127:112]),
.op_dout(op_dout_38_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_39_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_39[15:0]),
.op_dout(op_dout_39_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_39_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_39[31:16]),
.op_dout(op_dout_39_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_39_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_39[47:32]),
.op_dout(op_dout_39_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_39_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_39[63:48]),
.op_dout(op_dout_39_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_39_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_39[79:64]),
.op_dout(op_dout_39_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_39_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_39[95:80]),
.op_dout(op_dout_39_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_39_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_39[111:96]),
.op_dout(op_dout_39_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_39_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_39[127:112]),
.op_dout(op_dout_39_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_40_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_40[15:0]),
.op_dout(op_dout_40_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_40_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_40[31:16]),
.op_dout(op_dout_40_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_40_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_40[47:32]),
.op_dout(op_dout_40_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_40_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_40[63:48]),
.op_dout(op_dout_40_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_40_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_40[79:64]),
.op_dout(op_dout_40_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_40_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_40[95:80]),
.op_dout(op_dout_40_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_40_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_40[111:96]),
.op_dout(op_dout_40_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_40_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_40[127:112]),
.op_dout(op_dout_40_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_41_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_41[15:0]),
.op_dout(op_dout_41_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_41_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_41[31:16]),
.op_dout(op_dout_41_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_41_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_41[47:32]),
.op_dout(op_dout_41_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_41_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_41[63:48]),
.op_dout(op_dout_41_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_41_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_41[79:64]),
.op_dout(op_dout_41_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_41_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_41[95:80]),
.op_dout(op_dout_41_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_41_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_41[111:96]),
.op_dout(op_dout_41_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_41_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_41[127:112]),
.op_dout(op_dout_41_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_42_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_42[15:0]),
.op_dout(op_dout_42_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_42_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_42[31:16]),
.op_dout(op_dout_42_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_42_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_42[47:32]),
.op_dout(op_dout_42_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_42_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_42[63:48]),
.op_dout(op_dout_42_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_42_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_42[79:64]),
.op_dout(op_dout_42_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_42_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_42[95:80]),
.op_dout(op_dout_42_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_42_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_42[111:96]),
.op_dout(op_dout_42_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_42_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_42[127:112]),
.op_dout(op_dout_42_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_43_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_43[15:0]),
.op_dout(op_dout_43_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_43_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_43[31:16]),
.op_dout(op_dout_43_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_43_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_43[47:32]),
.op_dout(op_dout_43_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_43_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_43[63:48]),
.op_dout(op_dout_43_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_43_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_43[79:64]),
.op_dout(op_dout_43_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_43_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_43[95:80]),
.op_dout(op_dout_43_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_43_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_43[111:96]),
.op_dout(op_dout_43_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_43_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_43[127:112]),
.op_dout(op_dout_43_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_44_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_44[15:0]),
.op_dout(op_dout_44_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_44_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_44[31:16]),
.op_dout(op_dout_44_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_44_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_44[47:32]),
.op_dout(op_dout_44_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_44_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_44[63:48]),
.op_dout(op_dout_44_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_44_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_44[79:64]),
.op_dout(op_dout_44_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_44_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_44[95:80]),
.op_dout(op_dout_44_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_44_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_44[111:96]),
.op_dout(op_dout_44_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_44_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_44[127:112]),
.op_dout(op_dout_44_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_45_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_45[15:0]),
.op_dout(op_dout_45_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_45_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_45[31:16]),
.op_dout(op_dout_45_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_45_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_45[47:32]),
.op_dout(op_dout_45_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_45_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_45[63:48]),
.op_dout(op_dout_45_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_45_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_45[79:64]),
.op_dout(op_dout_45_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_45_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_45[95:80]),
.op_dout(op_dout_45_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_45_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_45[111:96]),
.op_dout(op_dout_45_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_45_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_45[127:112]),
.op_dout(op_dout_45_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_46_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_46[15:0]),
.op_dout(op_dout_46_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_46_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_46[31:16]),
.op_dout(op_dout_46_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_46_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_46[47:32]),
.op_dout(op_dout_46_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_46_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_46[63:48]),
.op_dout(op_dout_46_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_46_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_46[79:64]),
.op_dout(op_dout_46_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_46_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_46[95:80]),
.op_dout(op_dout_46_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_46_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_46[111:96]),
.op_dout(op_dout_46_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_46_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_46[127:112]),
.op_dout(op_dout_46_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_47_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_47[15:0]),
.op_dout(op_dout_47_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_47_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_47[31:16]),
.op_dout(op_dout_47_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_47_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_47[47:32]),
.op_dout(op_dout_47_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_47_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_47[63:48]),
.op_dout(op_dout_47_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_47_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_47[79:64]),
.op_dout(op_dout_47_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_47_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_47[95:80]),
.op_dout(op_dout_47_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_47_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_47[111:96]),
.op_dout(op_dout_47_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_47_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_47[127:112]),
.op_dout(op_dout_47_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_48_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_48[15:0]),
.op_dout(op_dout_48_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_48_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_48[31:16]),
.op_dout(op_dout_48_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_48_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_48[47:32]),
.op_dout(op_dout_48_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_48_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_48[63:48]),
.op_dout(op_dout_48_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_48_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_48[79:64]),
.op_dout(op_dout_48_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_48_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_48[95:80]),
.op_dout(op_dout_48_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_48_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_48[111:96]),
.op_dout(op_dout_48_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_48_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_48[127:112]),
.op_dout(op_dout_48_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_49_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_49[15:0]),
.op_dout(op_dout_49_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_49_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_49[31:16]),
.op_dout(op_dout_49_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_49_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_49[47:32]),
.op_dout(op_dout_49_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_49_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_49[63:48]),
.op_dout(op_dout_49_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_49_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_49[79:64]),
.op_dout(op_dout_49_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_49_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_49[95:80]),
.op_dout(op_dout_49_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_49_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_49[111:96]),
.op_dout(op_dout_49_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_49_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_49[127:112]),
.op_dout(op_dout_49_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_50_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_50[15:0]),
.op_dout(op_dout_50_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_50_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_50[31:16]),
.op_dout(op_dout_50_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_50_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_50[47:32]),
.op_dout(op_dout_50_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_50_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_50[63:48]),
.op_dout(op_dout_50_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_50_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_50[79:64]),
.op_dout(op_dout_50_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_50_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_50[95:80]),
.op_dout(op_dout_50_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_50_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_50[111:96]),
.op_dout(op_dout_50_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_50_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_50[127:112]),
.op_dout(op_dout_50_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_51_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_51[15:0]),
.op_dout(op_dout_51_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_51_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_51[31:16]),
.op_dout(op_dout_51_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_51_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_51[47:32]),
.op_dout(op_dout_51_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_51_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_51[63:48]),
.op_dout(op_dout_51_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_51_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_51[79:64]),
.op_dout(op_dout_51_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_51_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_51[95:80]),
.op_dout(op_dout_51_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_51_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_51[111:96]),
.op_dout(op_dout_51_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_51_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_51[127:112]),
.op_dout(op_dout_51_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_52_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_52[15:0]),
.op_dout(op_dout_52_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_52_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_52[31:16]),
.op_dout(op_dout_52_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_52_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_52[47:32]),
.op_dout(op_dout_52_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_52_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_52[63:48]),
.op_dout(op_dout_52_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_52_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_52[79:64]),
.op_dout(op_dout_52_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_52_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_52[95:80]),
.op_dout(op_dout_52_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_52_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_52[111:96]),
.op_dout(op_dout_52_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_52_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_52[127:112]),
.op_dout(op_dout_52_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_53_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_53[15:0]),
.op_dout(op_dout_53_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_53_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_53[31:16]),
.op_dout(op_dout_53_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_53_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_53[47:32]),
.op_dout(op_dout_53_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_53_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_53[63:48]),
.op_dout(op_dout_53_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_53_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_53[79:64]),
.op_dout(op_dout_53_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_53_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_53[95:80]),
.op_dout(op_dout_53_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_53_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_53[111:96]),
.op_dout(op_dout_53_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_53_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_53[127:112]),
.op_dout(op_dout_53_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_54_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_54[15:0]),
.op_dout(op_dout_54_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_54_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_54[31:16]),
.op_dout(op_dout_54_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_54_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_54[47:32]),
.op_dout(op_dout_54_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_54_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_54[63:48]),
.op_dout(op_dout_54_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_54_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_54[79:64]),
.op_dout(op_dout_54_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_54_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_54[95:80]),
.op_dout(op_dout_54_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_54_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_54[111:96]),
.op_dout(op_dout_54_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_54_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_54[127:112]),
.op_dout(op_dout_54_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_55_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_55[15:0]),
.op_dout(op_dout_55_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_55_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_55[31:16]),
.op_dout(op_dout_55_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_55_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_55[47:32]),
.op_dout(op_dout_55_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_55_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_55[63:48]),
.op_dout(op_dout_55_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_55_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_55[79:64]),
.op_dout(op_dout_55_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_55_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_55[95:80]),
.op_dout(op_dout_55_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_55_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_55[111:96]),
.op_dout(op_dout_55_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_55_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_55[127:112]),
.op_dout(op_dout_55_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_56_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_56[15:0]),
.op_dout(op_dout_56_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_56_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_56[31:16]),
.op_dout(op_dout_56_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_56_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_56[47:32]),
.op_dout(op_dout_56_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_56_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_56[63:48]),
.op_dout(op_dout_56_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_56_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_56[79:64]),
.op_dout(op_dout_56_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_56_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_56[95:80]),
.op_dout(op_dout_56_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_56_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_56[111:96]),
.op_dout(op_dout_56_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_56_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_56[127:112]),
.op_dout(op_dout_56_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_57_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_57[15:0]),
.op_dout(op_dout_57_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_57_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_57[31:16]),
.op_dout(op_dout_57_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_57_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_57[47:32]),
.op_dout(op_dout_57_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_57_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_57[63:48]),
.op_dout(op_dout_57_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_57_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_57[79:64]),
.op_dout(op_dout_57_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_57_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_57[95:80]),
.op_dout(op_dout_57_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_57_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_57[111:96]),
.op_dout(op_dout_57_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_57_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_57[127:112]),
.op_dout(op_dout_57_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_58_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_58[15:0]),
.op_dout(op_dout_58_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_58_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_58[31:16]),
.op_dout(op_dout_58_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_58_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_58[47:32]),
.op_dout(op_dout_58_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_58_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_58[63:48]),
.op_dout(op_dout_58_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_58_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_58[79:64]),
.op_dout(op_dout_58_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_58_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_58[95:80]),
.op_dout(op_dout_58_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_58_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_58[111:96]),
.op_dout(op_dout_58_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_58_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_58[127:112]),
.op_dout(op_dout_58_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_59_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_59[15:0]),
.op_dout(op_dout_59_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_59_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_59[31:16]),
.op_dout(op_dout_59_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_59_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_59[47:32]),
.op_dout(op_dout_59_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_59_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_59[63:48]),
.op_dout(op_dout_59_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_59_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_59[79:64]),
.op_dout(op_dout_59_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_59_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_59[95:80]),
.op_dout(op_dout_59_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_59_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_59[111:96]),
.op_dout(op_dout_59_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_59_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_59[127:112]),
.op_dout(op_dout_59_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_60_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_60[15:0]),
.op_dout(op_dout_60_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_60_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_60[31:16]),
.op_dout(op_dout_60_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_60_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_60[47:32]),
.op_dout(op_dout_60_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_60_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_60[63:48]),
.op_dout(op_dout_60_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_60_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_60[79:64]),
.op_dout(op_dout_60_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_60_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_60[95:80]),
.op_dout(op_dout_60_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_60_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_60[111:96]),
.op_dout(op_dout_60_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_60_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_60[127:112]),
.op_dout(op_dout_60_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_61_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_61[15:0]),
.op_dout(op_dout_61_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_61_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_61[31:16]),
.op_dout(op_dout_61_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_61_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_61[47:32]),
.op_dout(op_dout_61_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_61_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_61[63:48]),
.op_dout(op_dout_61_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_61_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_61[79:64]),
.op_dout(op_dout_61_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_61_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_61[95:80]),
.op_dout(op_dout_61_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_61_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_61[111:96]),
.op_dout(op_dout_61_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_61_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_61[127:112]),
.op_dout(op_dout_61_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_62_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_62[15:0]),
.op_dout(op_dout_62_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_62_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_62[31:16]),
.op_dout(op_dout_62_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_62_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_62[47:32]),
.op_dout(op_dout_62_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_62_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_62[63:48]),
.op_dout(op_dout_62_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_62_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_62[79:64]),
.op_dout(op_dout_62_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_62_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_62[95:80]),
.op_dout(op_dout_62_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_62_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_62[111:96]),
.op_dout(op_dout_62_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_62_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_62[127:112]),
.op_dout(op_dout_62_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_63_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_63[15:0]),
.op_dout(op_dout_63_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_63_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_63[31:16]),
.op_dout(op_dout_63_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_63_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_63[47:32]),
.op_dout(op_dout_63_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_63_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_63[63:48]),
.op_dout(op_dout_63_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_63_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_63[79:64]),
.op_dout(op_dout_63_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_63_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_63[95:80]),
.op_dout(op_dout_63_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_63_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_63[111:96]),
.op_dout(op_dout_63_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_63_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_63[127:112]),
.op_dout(op_dout_63_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_64_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_64[15:0]),
.op_dout(op_dout_64_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_64_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_64[31:16]),
.op_dout(op_dout_64_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_64_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_64[47:32]),
.op_dout(op_dout_64_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_64_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_64[63:48]),
.op_dout(op_dout_64_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_64_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_64[79:64]),
.op_dout(op_dout_64_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_64_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_64[95:80]),
.op_dout(op_dout_64_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_64_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_64[111:96]),
.op_dout(op_dout_64_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_64_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_64[127:112]),
.op_dout(op_dout_64_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_65_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_65[15:0]),
.op_dout(op_dout_65_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_65_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_65[31:16]),
.op_dout(op_dout_65_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_65_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_65[47:32]),
.op_dout(op_dout_65_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_65_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_65[63:48]),
.op_dout(op_dout_65_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_65_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_65[79:64]),
.op_dout(op_dout_65_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_65_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_65[95:80]),
.op_dout(op_dout_65_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_65_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_65[111:96]),
.op_dout(op_dout_65_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_65_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_65[127:112]),
.op_dout(op_dout_65_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_66_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_66[15:0]),
.op_dout(op_dout_66_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_66_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_66[31:16]),
.op_dout(op_dout_66_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_66_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_66[47:32]),
.op_dout(op_dout_66_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_66_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_66[63:48]),
.op_dout(op_dout_66_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_66_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_66[79:64]),
.op_dout(op_dout_66_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_66_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_66[95:80]),
.op_dout(op_dout_66_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_66_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_66[111:96]),
.op_dout(op_dout_66_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_66_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_66[127:112]),
.op_dout(op_dout_66_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_67_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_67[15:0]),
.op_dout(op_dout_67_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_67_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_67[31:16]),
.op_dout(op_dout_67_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_67_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_67[47:32]),
.op_dout(op_dout_67_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_67_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_67[63:48]),
.op_dout(op_dout_67_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_67_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_67[79:64]),
.op_dout(op_dout_67_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_67_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_67[95:80]),
.op_dout(op_dout_67_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_67_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_67[111:96]),
.op_dout(op_dout_67_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_67_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_67[127:112]),
.op_dout(op_dout_67_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_68_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_68[15:0]),
.op_dout(op_dout_68_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_68_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_68[31:16]),
.op_dout(op_dout_68_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_68_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_68[47:32]),
.op_dout(op_dout_68_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_68_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_68[63:48]),
.op_dout(op_dout_68_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_68_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_68[79:64]),
.op_dout(op_dout_68_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_68_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_68[95:80]),
.op_dout(op_dout_68_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_68_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_68[111:96]),
.op_dout(op_dout_68_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_68_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_68[127:112]),
.op_dout(op_dout_68_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_69_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_69[15:0]),
.op_dout(op_dout_69_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_69_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_69[31:16]),
.op_dout(op_dout_69_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_69_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_69[47:32]),
.op_dout(op_dout_69_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_69_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_69[63:48]),
.op_dout(op_dout_69_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_69_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_69[79:64]),
.op_dout(op_dout_69_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_69_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_69[95:80]),
.op_dout(op_dout_69_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_69_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_69[111:96]),
.op_dout(op_dout_69_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_69_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_69[127:112]),
.op_dout(op_dout_69_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_70_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_70[15:0]),
.op_dout(op_dout_70_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_70_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_70[31:16]),
.op_dout(op_dout_70_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_70_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_70[47:32]),
.op_dout(op_dout_70_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_70_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_70[63:48]),
.op_dout(op_dout_70_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_70_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_70[79:64]),
.op_dout(op_dout_70_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_70_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_70[95:80]),
.op_dout(op_dout_70_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_70_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_70[111:96]),
.op_dout(op_dout_70_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_70_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_70[127:112]),
.op_dout(op_dout_70_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_71_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_71[15:0]),
.op_dout(op_dout_71_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_71_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_71[31:16]),
.op_dout(op_dout_71_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_71_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_71[47:32]),
.op_dout(op_dout_71_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_71_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_71[63:48]),
.op_dout(op_dout_71_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_71_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_71[79:64]),
.op_dout(op_dout_71_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_71_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_71[95:80]),
.op_dout(op_dout_71_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_71_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_71[111:96]),
.op_dout(op_dout_71_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_71_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_71[127:112]),
.op_dout(op_dout_71_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_72_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_72[15:0]),
.op_dout(op_dout_72_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_72_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_72[31:16]),
.op_dout(op_dout_72_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_72_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_72[47:32]),
.op_dout(op_dout_72_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_72_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_72[63:48]),
.op_dout(op_dout_72_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_72_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_72[79:64]),
.op_dout(op_dout_72_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_72_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_72[95:80]),
.op_dout(op_dout_72_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_72_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_72[111:96]),
.op_dout(op_dout_72_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_72_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_72[127:112]),
.op_dout(op_dout_72_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_73_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_73[15:0]),
.op_dout(op_dout_73_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_73_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_73[31:16]),
.op_dout(op_dout_73_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_73_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_73[47:32]),
.op_dout(op_dout_73_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_73_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_73[63:48]),
.op_dout(op_dout_73_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_73_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_73[79:64]),
.op_dout(op_dout_73_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_73_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_73[95:80]),
.op_dout(op_dout_73_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_73_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_73[111:96]),
.op_dout(op_dout_73_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_73_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_73[127:112]),
.op_dout(op_dout_73_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_74_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_74[15:0]),
.op_dout(op_dout_74_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_74_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_74[31:16]),
.op_dout(op_dout_74_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_74_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_74[47:32]),
.op_dout(op_dout_74_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_74_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_74[63:48]),
.op_dout(op_dout_74_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_74_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_74[79:64]),
.op_dout(op_dout_74_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_74_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_74[95:80]),
.op_dout(op_dout_74_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_74_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_74[111:96]),
.op_dout(op_dout_74_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_74_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_74[127:112]),
.op_dout(op_dout_74_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_75_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_75[15:0]),
.op_dout(op_dout_75_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_75_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_75[31:16]),
.op_dout(op_dout_75_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_75_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_75[47:32]),
.op_dout(op_dout_75_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_75_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_75[63:48]),
.op_dout(op_dout_75_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_75_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_75[79:64]),
.op_dout(op_dout_75_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_75_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_75[95:80]),
.op_dout(op_dout_75_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_75_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_75[111:96]),
.op_dout(op_dout_75_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_75_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_75[127:112]),
.op_dout(op_dout_75_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_76_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_76[15:0]),
.op_dout(op_dout_76_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_76_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_76[31:16]),
.op_dout(op_dout_76_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_76_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_76[47:32]),
.op_dout(op_dout_76_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_76_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_76[63:48]),
.op_dout(op_dout_76_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_76_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_76[79:64]),
.op_dout(op_dout_76_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_76_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_76[95:80]),
.op_dout(op_dout_76_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_76_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_76[111:96]),
.op_dout(op_dout_76_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_76_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_76[127:112]),
.op_dout(op_dout_76_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_77_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_77[15:0]),
.op_dout(op_dout_77_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_77_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_77[31:16]),
.op_dout(op_dout_77_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_77_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_77[47:32]),
.op_dout(op_dout_77_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_77_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_77[63:48]),
.op_dout(op_dout_77_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_77_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_77[79:64]),
.op_dout(op_dout_77_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_77_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_77[95:80]),
.op_dout(op_dout_77_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_77_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_77[111:96]),
.op_dout(op_dout_77_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_77_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_77[127:112]),
.op_dout(op_dout_77_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_78_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_78[15:0]),
.op_dout(op_dout_78_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_78_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_78[31:16]),
.op_dout(op_dout_78_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_78_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_78[47:32]),
.op_dout(op_dout_78_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_78_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_78[63:48]),
.op_dout(op_dout_78_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_78_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_78[79:64]),
.op_dout(op_dout_78_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_78_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_78[95:80]),
.op_dout(op_dout_78_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_78_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_78[111:96]),
.op_dout(op_dout_78_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_78_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_78[127:112]),
.op_dout(op_dout_78_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_79_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_79[15:0]),
.op_dout(op_dout_79_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_79_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_79[31:16]),
.op_dout(op_dout_79_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_79_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_79[47:32]),
.op_dout(op_dout_79_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_79_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_79[63:48]),
.op_dout(op_dout_79_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_79_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_79[79:64]),
.op_dout(op_dout_79_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_79_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_79[95:80]),
.op_dout(op_dout_79_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_79_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_79[111:96]),
.op_dout(op_dout_79_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_79_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_79[127:112]),
.op_dout(op_dout_79_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_80_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_80[15:0]),
.op_dout(op_dout_80_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_80_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_80[31:16]),
.op_dout(op_dout_80_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_80_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_80[47:32]),
.op_dout(op_dout_80_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_80_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_80[63:48]),
.op_dout(op_dout_80_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_80_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_80[79:64]),
.op_dout(op_dout_80_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_80_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_80[95:80]),
.op_dout(op_dout_80_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_80_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_80[111:96]),
.op_dout(op_dout_80_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_80_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_80[127:112]),
.op_dout(op_dout_80_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_81_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_81[15:0]),
.op_dout(op_dout_81_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_81_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_81[31:16]),
.op_dout(op_dout_81_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_81_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_81[47:32]),
.op_dout(op_dout_81_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_81_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_81[63:48]),
.op_dout(op_dout_81_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_81_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_81[79:64]),
.op_dout(op_dout_81_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_81_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_81[95:80]),
.op_dout(op_dout_81_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_81_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_81[111:96]),
.op_dout(op_dout_81_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_81_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_81[127:112]),
.op_dout(op_dout_81_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_82_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_82[15:0]),
.op_dout(op_dout_82_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_82_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_82[31:16]),
.op_dout(op_dout_82_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_82_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_82[47:32]),
.op_dout(op_dout_82_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_82_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_82[63:48]),
.op_dout(op_dout_82_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_82_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_82[79:64]),
.op_dout(op_dout_82_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_82_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_82[95:80]),
.op_dout(op_dout_82_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_82_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_82[111:96]),
.op_dout(op_dout_82_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_82_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_82[127:112]),
.op_dout(op_dout_82_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_83_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_83[15:0]),
.op_dout(op_dout_83_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_83_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_83[31:16]),
.op_dout(op_dout_83_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_83_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_83[47:32]),
.op_dout(op_dout_83_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_83_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_83[63:48]),
.op_dout(op_dout_83_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_83_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_83[79:64]),
.op_dout(op_dout_83_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_83_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_83[95:80]),
.op_dout(op_dout_83_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_83_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_83[111:96]),
.op_dout(op_dout_83_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_83_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_83[127:112]),
.op_dout(op_dout_83_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_84_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_84[15:0]),
.op_dout(op_dout_84_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_84_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_84[31:16]),
.op_dout(op_dout_84_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_84_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_84[47:32]),
.op_dout(op_dout_84_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_84_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_84[63:48]),
.op_dout(op_dout_84_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_84_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_84[79:64]),
.op_dout(op_dout_84_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_84_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_84[95:80]),
.op_dout(op_dout_84_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_84_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_84[111:96]),
.op_dout(op_dout_84_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_84_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_84[127:112]),
.op_dout(op_dout_84_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_85_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_85[15:0]),
.op_dout(op_dout_85_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_85_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_85[31:16]),
.op_dout(op_dout_85_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_85_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_85[47:32]),
.op_dout(op_dout_85_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_85_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_85[63:48]),
.op_dout(op_dout_85_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_85_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_85[79:64]),
.op_dout(op_dout_85_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_85_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_85[95:80]),
.op_dout(op_dout_85_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_85_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_85[111:96]),
.op_dout(op_dout_85_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_85_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_85[127:112]),
.op_dout(op_dout_85_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_86_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_86[15:0]),
.op_dout(op_dout_86_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_86_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_86[31:16]),
.op_dout(op_dout_86_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_86_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_86[47:32]),
.op_dout(op_dout_86_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_86_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_86[63:48]),
.op_dout(op_dout_86_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_86_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_86[79:64]),
.op_dout(op_dout_86_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_86_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_86[95:80]),
.op_dout(op_dout_86_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_86_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_86[111:96]),
.op_dout(op_dout_86_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_86_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_86[127:112]),
.op_dout(op_dout_86_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_87_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_87[15:0]),
.op_dout(op_dout_87_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_87_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_87[31:16]),
.op_dout(op_dout_87_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_87_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_87[47:32]),
.op_dout(op_dout_87_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_87_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_87[63:48]),
.op_dout(op_dout_87_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_87_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_87[79:64]),
.op_dout(op_dout_87_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_87_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_87[95:80]),
.op_dout(op_dout_87_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_87_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_87[111:96]),
.op_dout(op_dout_87_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_87_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_87[127:112]),
.op_dout(op_dout_87_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_88_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_88[15:0]),
.op_dout(op_dout_88_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_88_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_88[31:16]),
.op_dout(op_dout_88_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_88_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_88[47:32]),
.op_dout(op_dout_88_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_88_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_88[63:48]),
.op_dout(op_dout_88_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_88_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_88[79:64]),
.op_dout(op_dout_88_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_88_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_88[95:80]),
.op_dout(op_dout_88_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_88_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_88[111:96]),
.op_dout(op_dout_88_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_88_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_88[127:112]),
.op_dout(op_dout_88_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_89_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_89[15:0]),
.op_dout(op_dout_89_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_89_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_89[31:16]),
.op_dout(op_dout_89_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_89_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_89[47:32]),
.op_dout(op_dout_89_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_89_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_89[63:48]),
.op_dout(op_dout_89_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_89_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_89[79:64]),
.op_dout(op_dout_89_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_89_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_89[95:80]),
.op_dout(op_dout_89_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_89_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_89[111:96]),
.op_dout(op_dout_89_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_89_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_89[127:112]),
.op_dout(op_dout_89_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_90_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_90[15:0]),
.op_dout(op_dout_90_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_90_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_90[31:16]),
.op_dout(op_dout_90_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_90_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_90[47:32]),
.op_dout(op_dout_90_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_90_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_90[63:48]),
.op_dout(op_dout_90_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_90_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_90[79:64]),
.op_dout(op_dout_90_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_90_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_90[95:80]),
.op_dout(op_dout_90_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_90_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_90[111:96]),
.op_dout(op_dout_90_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_90_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_90[127:112]),
.op_dout(op_dout_90_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_91_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_91[15:0]),
.op_dout(op_dout_91_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_91_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_91[31:16]),
.op_dout(op_dout_91_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_91_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_91[47:32]),
.op_dout(op_dout_91_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_91_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_91[63:48]),
.op_dout(op_dout_91_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_91_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_91[79:64]),
.op_dout(op_dout_91_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_91_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_91[95:80]),
.op_dout(op_dout_91_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_91_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_91[111:96]),
.op_dout(op_dout_91_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_91_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_91[127:112]),
.op_dout(op_dout_91_7));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_92_0(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_92[15:0]),
.op_dout(op_dout_92_0));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_92_1(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_92[31:16]),
.op_dout(op_dout_92_1));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_92_2(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_92[47:32]),
.op_dout(op_dout_92_2));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_92_3(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_92[63:48]),
.op_dout(op_dout_92_3));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_92_4(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_92[79:64]),
.op_dout(op_dout_92_4));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_92_5(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_92[95:80]),
.op_dout(op_dout_92_5));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_92_6(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_92[111:96]),
.op_dout(op_dout_92_6));

vector_max #(.RELU(0),
.DIN_W(16),
.Q(13))
u_vector_max_92_7(
.clk(clk),
.rst(rst),
.op_din_en(op_din_en),
.op_din_eop(op_din_eop),
.op_din(op_data_92[127:112]),
.op_dout(op_dout_92_7));

assign blob_dout_fifo = {op_dout_92_7,op_dout_92_6,op_dout_92_5,op_dout_92_4,op_dout_92_3,op_dout_92_2,op_dout_92_1,op_dout_92_0,op_dout_91_7,op_dout_91_6,op_dout_91_5,op_dout_91_4,op_dout_91_3,op_dout_91_2,op_dout_91_1,op_dout_91_0,op_dout_90_7,op_dout_90_6,op_dout_90_5,op_dout_90_4,op_dout_90_3,op_dout_90_2,op_dout_90_1,op_dout_90_0,op_dout_89_7,op_dout_89_6,op_dout_89_5,op_dout_89_4,op_dout_89_3,op_dout_89_2,op_dout_89_1,op_dout_89_0,op_dout_88_7,op_dout_88_6,op_dout_88_5,op_dout_88_4,op_dout_88_3,op_dout_88_2,op_dout_88_1,op_dout_88_0,op_dout_87_7,op_dout_87_6,op_dout_87_5,op_dout_87_4,op_dout_87_3,op_dout_87_2,op_dout_87_1,op_dout_87_0,op_dout_86_7,op_dout_86_6,op_dout_86_5,op_dout_86_4,op_dout_86_3,op_dout_86_2,op_dout_86_1,op_dout_86_0,op_dout_85_7,op_dout_85_6,op_dout_85_5,op_dout_85_4,op_dout_85_3,op_dout_85_2,op_dout_85_1,op_dout_85_0,op_dout_84_7,op_dout_84_6,op_dout_84_5,op_dout_84_4,op_dout_84_3,op_dout_84_2,op_dout_84_1,op_dout_84_0,op_dout_83_7,op_dout_83_6,op_dout_83_5,op_dout_83_4,op_dout_83_3,op_dout_83_2,op_dout_83_1,op_dout_83_0,op_dout_82_7,op_dout_82_6,op_dout_82_5,op_dout_82_4,op_dout_82_3,op_dout_82_2,op_dout_82_1,op_dout_82_0,op_dout_81_7,op_dout_81_6,op_dout_81_5,op_dout_81_4,op_dout_81_3,op_dout_81_2,op_dout_81_1,op_dout_81_0,op_dout_80_7,op_dout_80_6,op_dout_80_5,op_dout_80_4,op_dout_80_3,op_dout_80_2,op_dout_80_1,op_dout_80_0,op_dout_79_7,op_dout_79_6,op_dout_79_5,op_dout_79_4,op_dout_79_3,op_dout_79_2,op_dout_79_1,op_dout_79_0,op_dout_78_7,op_dout_78_6,op_dout_78_5,op_dout_78_4,op_dout_78_3,op_dout_78_2,op_dout_78_1,op_dout_78_0,op_dout_77_7,op_dout_77_6,op_dout_77_5,op_dout_77_4,op_dout_77_3,op_dout_77_2,op_dout_77_1,op_dout_77_0,op_dout_76_7,op_dout_76_6,op_dout_76_5,op_dout_76_4,op_dout_76_3,op_dout_76_2,op_dout_76_1,op_dout_76_0,op_dout_75_7,op_dout_75_6,op_dout_75_5,op_dout_75_4,op_dout_75_3,op_dout_75_2,op_dout_75_1,op_dout_75_0,op_dout_74_7,op_dout_74_6,op_dout_74_5,op_dout_74_4,op_dout_74_3,op_dout_74_2,op_dout_74_1,op_dout_74_0,op_dout_73_7,op_dout_73_6,op_dout_73_5,op_dout_73_4,op_dout_73_3,op_dout_73_2,op_dout_73_1,op_dout_73_0,op_dout_72_7,op_dout_72_6,op_dout_72_5,op_dout_72_4,op_dout_72_3,op_dout_72_2,op_dout_72_1,op_dout_72_0,op_dout_71_7,op_dout_71_6,op_dout_71_5,op_dout_71_4,op_dout_71_3,op_dout_71_2,op_dout_71_1,op_dout_71_0,op_dout_70_7,op_dout_70_6,op_dout_70_5,op_dout_70_4,op_dout_70_3,op_dout_70_2,op_dout_70_1,op_dout_70_0,op_dout_69_7,op_dout_69_6,op_dout_69_5,op_dout_69_4,op_dout_69_3,op_dout_69_2,op_dout_69_1,op_dout_69_0,op_dout_68_7,op_dout_68_6,op_dout_68_5,op_dout_68_4,op_dout_68_3,op_dout_68_2,op_dout_68_1,op_dout_68_0,op_dout_67_7,op_dout_67_6,op_dout_67_5,op_dout_67_4,op_dout_67_3,op_dout_67_2,op_dout_67_1,op_dout_67_0,op_dout_66_7,op_dout_66_6,op_dout_66_5,op_dout_66_4,op_dout_66_3,op_dout_66_2,op_dout_66_1,op_dout_66_0,op_dout_65_7,op_dout_65_6,op_dout_65_5,op_dout_65_4,op_dout_65_3,op_dout_65_2,op_dout_65_1,op_dout_65_0,op_dout_64_7,op_dout_64_6,op_dout_64_5,op_dout_64_4,op_dout_64_3,op_dout_64_2,op_dout_64_1,op_dout_64_0,op_dout_63_7,op_dout_63_6,op_dout_63_5,op_dout_63_4,op_dout_63_3,op_dout_63_2,op_dout_63_1,op_dout_63_0,op_dout_62_7,op_dout_62_6,op_dout_62_5,op_dout_62_4,op_dout_62_3,op_dout_62_2,op_dout_62_1,op_dout_62_0,op_dout_61_7,op_dout_61_6,op_dout_61_5,op_dout_61_4,op_dout_61_3,op_dout_61_2,op_dout_61_1,op_dout_61_0,op_dout_60_7,op_dout_60_6,op_dout_60_5,op_dout_60_4,op_dout_60_3,op_dout_60_2,op_dout_60_1,op_dout_60_0,op_dout_59_7,op_dout_59_6,op_dout_59_5,op_dout_59_4,op_dout_59_3,op_dout_59_2,op_dout_59_1,op_dout_59_0,op_dout_58_7,op_dout_58_6,op_dout_58_5,op_dout_58_4,op_dout_58_3,op_dout_58_2,op_dout_58_1,op_dout_58_0,op_dout_57_7,op_dout_57_6,op_dout_57_5,op_dout_57_4,op_dout_57_3,op_dout_57_2,op_dout_57_1,op_dout_57_0,op_dout_56_7,op_dout_56_6,op_dout_56_5,op_dout_56_4,op_dout_56_3,op_dout_56_2,op_dout_56_1,op_dout_56_0,op_dout_55_7,op_dout_55_6,op_dout_55_5,op_dout_55_4,op_dout_55_3,op_dout_55_2,op_dout_55_1,op_dout_55_0,op_dout_54_7,op_dout_54_6,op_dout_54_5,op_dout_54_4,op_dout_54_3,op_dout_54_2,op_dout_54_1,op_dout_54_0,op_dout_53_7,op_dout_53_6,op_dout_53_5,op_dout_53_4,op_dout_53_3,op_dout_53_2,op_dout_53_1,op_dout_53_0,op_dout_52_7,op_dout_52_6,op_dout_52_5,op_dout_52_4,op_dout_52_3,op_dout_52_2,op_dout_52_1,op_dout_52_0,op_dout_51_7,op_dout_51_6,op_dout_51_5,op_dout_51_4,op_dout_51_3,op_dout_51_2,op_dout_51_1,op_dout_51_0,op_dout_50_7,op_dout_50_6,op_dout_50_5,op_dout_50_4,op_dout_50_3,op_dout_50_2,op_dout_50_1,op_dout_50_0,op_dout_49_7,op_dout_49_6,op_dout_49_5,op_dout_49_4,op_dout_49_3,op_dout_49_2,op_dout_49_1,op_dout_49_0,op_dout_48_7,op_dout_48_6,op_dout_48_5,op_dout_48_4,op_dout_48_3,op_dout_48_2,op_dout_48_1,op_dout_48_0,op_dout_47_7,op_dout_47_6,op_dout_47_5,op_dout_47_4,op_dout_47_3,op_dout_47_2,op_dout_47_1,op_dout_47_0,op_dout_46_7,op_dout_46_6,op_dout_46_5,op_dout_46_4,op_dout_46_3,op_dout_46_2,op_dout_46_1,op_dout_46_0,op_dout_45_7,op_dout_45_6,op_dout_45_5,op_dout_45_4,op_dout_45_3,op_dout_45_2,op_dout_45_1,op_dout_45_0,op_dout_44_7,op_dout_44_6,op_dout_44_5,op_dout_44_4,op_dout_44_3,op_dout_44_2,op_dout_44_1,op_dout_44_0,op_dout_43_7,op_dout_43_6,op_dout_43_5,op_dout_43_4,op_dout_43_3,op_dout_43_2,op_dout_43_1,op_dout_43_0,op_dout_42_7,op_dout_42_6,op_dout_42_5,op_dout_42_4,op_dout_42_3,op_dout_42_2,op_dout_42_1,op_dout_42_0,op_dout_41_7,op_dout_41_6,op_dout_41_5,op_dout_41_4,op_dout_41_3,op_dout_41_2,op_dout_41_1,op_dout_41_0,op_dout_40_7,op_dout_40_6,op_dout_40_5,op_dout_40_4,op_dout_40_3,op_dout_40_2,op_dout_40_1,op_dout_40_0,op_dout_39_7,op_dout_39_6,op_dout_39_5,op_dout_39_4,op_dout_39_3,op_dout_39_2,op_dout_39_1,op_dout_39_0,op_dout_38_7,op_dout_38_6,op_dout_38_5,op_dout_38_4,op_dout_38_3,op_dout_38_2,op_dout_38_1,op_dout_38_0,op_dout_37_7,op_dout_37_6,op_dout_37_5,op_dout_37_4,op_dout_37_3,op_dout_37_2,op_dout_37_1,op_dout_37_0,op_dout_36_7,op_dout_36_6,op_dout_36_5,op_dout_36_4,op_dout_36_3,op_dout_36_2,op_dout_36_1,op_dout_36_0,op_dout_35_7,op_dout_35_6,op_dout_35_5,op_dout_35_4,op_dout_35_3,op_dout_35_2,op_dout_35_1,op_dout_35_0,op_dout_34_7,op_dout_34_6,op_dout_34_5,op_dout_34_4,op_dout_34_3,op_dout_34_2,op_dout_34_1,op_dout_34_0,op_dout_33_7,op_dout_33_6,op_dout_33_5,op_dout_33_4,op_dout_33_3,op_dout_33_2,op_dout_33_1,op_dout_33_0,op_dout_32_7,op_dout_32_6,op_dout_32_5,op_dout_32_4,op_dout_32_3,op_dout_32_2,op_dout_32_1,op_dout_32_0,op_dout_31_7,op_dout_31_6,op_dout_31_5,op_dout_31_4,op_dout_31_3,op_dout_31_2,op_dout_31_1,op_dout_31_0,op_dout_30_7,op_dout_30_6,op_dout_30_5,op_dout_30_4,op_dout_30_3,op_dout_30_2,op_dout_30_1,op_dout_30_0,op_dout_29_7,op_dout_29_6,op_dout_29_5,op_dout_29_4,op_dout_29_3,op_dout_29_2,op_dout_29_1,op_dout_29_0,op_dout_28_7,op_dout_28_6,op_dout_28_5,op_dout_28_4,op_dout_28_3,op_dout_28_2,op_dout_28_1,op_dout_28_0,op_dout_27_7,op_dout_27_6,op_dout_27_5,op_dout_27_4,op_dout_27_3,op_dout_27_2,op_dout_27_1,op_dout_27_0,op_dout_26_7,op_dout_26_6,op_dout_26_5,op_dout_26_4,op_dout_26_3,op_dout_26_2,op_dout_26_1,op_dout_26_0,op_dout_25_7,op_dout_25_6,op_dout_25_5,op_dout_25_4,op_dout_25_3,op_dout_25_2,op_dout_25_1,op_dout_25_0,op_dout_24_7,op_dout_24_6,op_dout_24_5,op_dout_24_4,op_dout_24_3,op_dout_24_2,op_dout_24_1,op_dout_24_0,op_dout_23_7,op_dout_23_6,op_dout_23_5,op_dout_23_4,op_dout_23_3,op_dout_23_2,op_dout_23_1,op_dout_23_0,op_dout_22_7,op_dout_22_6,op_dout_22_5,op_dout_22_4,op_dout_22_3,op_dout_22_2,op_dout_22_1,op_dout_22_0,op_dout_21_7,op_dout_21_6,op_dout_21_5,op_dout_21_4,op_dout_21_3,op_dout_21_2,op_dout_21_1,op_dout_21_0,op_dout_20_7,op_dout_20_6,op_dout_20_5,op_dout_20_4,op_dout_20_3,op_dout_20_2,op_dout_20_1,op_dout_20_0,op_dout_19_7,op_dout_19_6,op_dout_19_5,op_dout_19_4,op_dout_19_3,op_dout_19_2,op_dout_19_1,op_dout_19_0,op_dout_18_7,op_dout_18_6,op_dout_18_5,op_dout_18_4,op_dout_18_3,op_dout_18_2,op_dout_18_1,op_dout_18_0,op_dout_17_7,op_dout_17_6,op_dout_17_5,op_dout_17_4,op_dout_17_3,op_dout_17_2,op_dout_17_1,op_dout_17_0,op_dout_16_7,op_dout_16_6,op_dout_16_5,op_dout_16_4,op_dout_16_3,op_dout_16_2,op_dout_16_1,op_dout_16_0,op_dout_15_7,op_dout_15_6,op_dout_15_5,op_dout_15_4,op_dout_15_3,op_dout_15_2,op_dout_15_1,op_dout_15_0,op_dout_14_7,op_dout_14_6,op_dout_14_5,op_dout_14_4,op_dout_14_3,op_dout_14_2,op_dout_14_1,op_dout_14_0,op_dout_13_7,op_dout_13_6,op_dout_13_5,op_dout_13_4,op_dout_13_3,op_dout_13_2,op_dout_13_1,op_dout_13_0,op_dout_12_7,op_dout_12_6,op_dout_12_5,op_dout_12_4,op_dout_12_3,op_dout_12_2,op_dout_12_1,op_dout_12_0,op_dout_11_7,op_dout_11_6,op_dout_11_5,op_dout_11_4,op_dout_11_3,op_dout_11_2,op_dout_11_1,op_dout_11_0,op_dout_10_7,op_dout_10_6,op_dout_10_5,op_dout_10_4,op_dout_10_3,op_dout_10_2,op_dout_10_1,op_dout_10_0,op_dout_9_7,op_dout_9_6,op_dout_9_5,op_dout_9_4,op_dout_9_3,op_dout_9_2,op_dout_9_1,op_dout_9_0,op_dout_8_7,op_dout_8_6,op_dout_8_5,op_dout_8_4,op_dout_8_3,op_dout_8_2,op_dout_8_1,op_dout_8_0,op_dout_7_7,op_dout_7_6,op_dout_7_5,op_dout_7_4,op_dout_7_3,op_dout_7_2,op_dout_7_1,op_dout_7_0,op_dout_6_7,op_dout_6_6,op_dout_6_5,op_dout_6_4,op_dout_6_3,op_dout_6_2,op_dout_6_1,op_dout_6_0,op_dout_5_7,op_dout_5_6,op_dout_5_5,op_dout_5_4,op_dout_5_3,op_dout_5_2,op_dout_5_1,op_dout_5_0,op_dout_4_7,op_dout_4_6,op_dout_4_5,op_dout_4_4,op_dout_4_3,op_dout_4_2,op_dout_4_1,op_dout_4_0,op_dout_3_7,op_dout_3_6,op_dout_3_5,op_dout_3_4,op_dout_3_3,op_dout_3_2,op_dout_3_1,op_dout_3_0,op_dout_2_7,op_dout_2_6,op_dout_2_5,op_dout_2_4,op_dout_2_3,op_dout_2_2,op_dout_2_1,op_dout_2_0,op_dout_1_7,op_dout_1_6,op_dout_1_5,op_dout_1_4,op_dout_1_3,op_dout_1_2,op_dout_1_1,op_dout_1_0,op_dout_0_7,op_dout_0_6,op_dout_0_5,op_dout_0_4,op_dout_0_3,op_dout_0_2,op_dout_0_1,op_dout_0_0};

wire empty_fifo;
wire blob_dout_eop_tmp;
assign blob_dout_en = blob_dout_rdy & (~empty_fifo);
assign blob_dout_eop = blob_dout_en & blob_dout_eop_tmp;
interlayer_sync_fifo #(
.aw(1),
.dw(11905),
.afull_t(2))
u_interlayer_sync_fifo (
.clk_i(clk),
.reset_i(rst),
.w_en_i(blob_dout_en_fifo), 
.w_din_i({blob_dout_eop_fifo, blob_dout_fifo}),
.r_en_i(blob_dout_en),
.r_dout_o({blob_dout_eop_tmp, blob_dout}),
.empty_o(empty_fifo),
.w_num_used_o(),
.r_num_val_o(),
.afull_o(),
.full_o());
endmodule
