VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO conv2_wm_sram_16_200_sky130A
   CLASS BLOCK ;
   SIZE 425.57 BY 357.74 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  128.52 0.0 129.26 1.93 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  141.61 0.0 142.35 1.93 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  155.89 0.0 156.63 1.93 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  168.98 0.0 169.72 1.93 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  182.07 0.0 182.81 1.93 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  193.97 0.0 194.71 1.93 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  208.25 0.0 208.99 1.93 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  221.34 0.0 222.08 1.93 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  234.43 0.0 235.17 1.93 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  247.52 0.0 248.26 1.93 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  260.61 0.0 261.35 1.93 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  273.7 0.0 274.44 1.93 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  286.79 0.0 287.53 1.93 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  299.88 0.0 300.62 1.93 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  312.97 0.0 313.71 1.93 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  327.25 0.0 327.99 1.93 ;
      END
   END din0[15]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  102.34 0.0 103.08 1.93 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  115.43 0.0 116.17 1.93 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 161.84 1.93 162.58 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 163.03 1.93 163.77 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 168.98 1.93 169.72 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 171.36 1.93 172.1 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 177.31 1.93 178.05 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 180.88 1.93 181.62 ;
      END
   END addr0[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 29.75 1.93 30.49 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 33.32 1.93 34.06 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  47.6 0.0 48.34 1.93 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  152.32 0.0 153.06 1.93 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  165.41 0.0 166.15 1.93 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  184.45 0.0 185.19 1.93 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  197.54 0.0 198.28 1.93 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  218.96 0.0 219.7 1.93 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  233.24 0.0 233.98 1.93 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  248.71 0.0 249.45 1.93 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  264.18 0.0 264.92 1.93 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  280.84 0.0 281.58 1.93 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  297.5 0.0 298.24 1.93 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  314.16 0.0 314.9 1.93 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  328.44 0.0 329.18 1.93 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  345.1 0.0 345.84 1.93 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  360.57 0.0 361.31 1.93 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  373.66 0.0 374.4 1.93 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  423.64 35.7 425.57 36.44 ;
      END
   END dout0[15]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  8.33 348.67 417.24 351.79 ;
         LAYER m4 ;
         RECT  8.33 8.33 11.45 351.79 ;
         LAYER m3 ;
         RECT  8.33 8.33 417.24 11.45 ;
         LAYER m4 ;
         RECT  414.12 8.33 417.24 351.79 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  2.38 2.38 423.19 5.5 ;
         LAYER m4 ;
         RECT  2.38 2.38 5.5 357.74 ;
         LAYER m4 ;
         RECT  420.07 2.38 423.19 357.74 ;
         LAYER m3 ;
         RECT  2.38 354.62 423.19 357.74 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  0.91 0.91 424.66 356.83 ;
   LAYER  m2 ;
      RECT  0.91 0.91 424.66 356.83 ;
   LAYER  m3 ;
      RECT  2.83 160.94 424.66 163.48 ;
      RECT  0.91 164.67 2.83 168.08 ;
      RECT  0.91 173.0 2.83 176.41 ;
      RECT  0.91 178.95 2.83 179.98 ;
      RECT  0.91 31.39 2.83 32.42 ;
      RECT  0.91 34.96 2.83 160.94 ;
      RECT  2.83 34.8 422.74 37.34 ;
      RECT  2.83 37.34 422.74 160.94 ;
      RECT  422.74 37.34 424.66 160.94 ;
      RECT  2.83 163.48 7.43 347.77 ;
      RECT  2.83 347.77 7.43 352.69 ;
      RECT  7.43 163.48 418.14 347.77 ;
      RECT  418.14 163.48 424.66 347.77 ;
      RECT  418.14 347.77 424.66 352.69 ;
      RECT  2.83 7.43 7.43 12.35 ;
      RECT  2.83 12.35 7.43 34.8 ;
      RECT  7.43 12.35 418.14 34.8 ;
      RECT  418.14 7.43 422.74 12.35 ;
      RECT  418.14 12.35 422.74 34.8 ;
      RECT  0.91 0.91 1.48 1.48 ;
      RECT  0.91 1.48 1.48 6.4 ;
      RECT  0.91 6.4 1.48 28.85 ;
      RECT  1.48 0.91 2.83 1.48 ;
      RECT  1.48 6.4 2.83 28.85 ;
      RECT  422.74 0.91 424.09 1.48 ;
      RECT  422.74 6.4 424.09 34.8 ;
      RECT  424.09 0.91 424.66 1.48 ;
      RECT  424.09 1.48 424.66 6.4 ;
      RECT  424.09 6.4 424.66 34.8 ;
      RECT  2.83 0.91 7.43 1.48 ;
      RECT  2.83 6.4 7.43 7.43 ;
      RECT  7.43 0.91 418.14 1.48 ;
      RECT  7.43 6.4 418.14 7.43 ;
      RECT  418.14 0.91 422.74 1.48 ;
      RECT  418.14 6.4 422.74 7.43 ;
      RECT  0.91 182.52 1.48 353.72 ;
      RECT  0.91 353.72 1.48 356.83 ;
      RECT  1.48 182.52 2.83 353.72 ;
      RECT  2.83 352.69 7.43 353.72 ;
      RECT  7.43 352.69 418.14 353.72 ;
      RECT  418.14 352.69 424.09 353.72 ;
      RECT  424.09 352.69 424.66 353.72 ;
      RECT  424.09 353.72 424.66 356.83 ;
   LAYER  m4 ;
      RECT  127.92 2.53 129.86 356.83 ;
      RECT  129.86 0.91 141.01 2.53 ;
      RECT  170.32 0.91 181.47 2.53 ;
      RECT  235.77 0.91 246.92 2.53 ;
      RECT  301.22 0.91 312.37 2.53 ;
      RECT  103.68 0.91 114.83 2.53 ;
      RECT  116.77 0.91 127.92 2.53 ;
      RECT  48.94 0.91 101.74 2.53 ;
      RECT  142.95 0.91 151.72 2.53 ;
      RECT  153.66 0.91 155.29 2.53 ;
      RECT  157.23 0.91 164.81 2.53 ;
      RECT  166.75 0.91 168.38 2.53 ;
      RECT  183.41 0.91 183.85 2.53 ;
      RECT  185.79 0.91 193.37 2.53 ;
      RECT  195.31 0.91 196.94 2.53 ;
      RECT  198.88 0.91 207.65 2.53 ;
      RECT  209.59 0.91 218.36 2.53 ;
      RECT  220.3 0.91 220.74 2.53 ;
      RECT  222.68 0.91 232.64 2.53 ;
      RECT  250.05 0.91 260.01 2.53 ;
      RECT  261.95 0.91 263.58 2.53 ;
      RECT  265.52 0.91 273.1 2.53 ;
      RECT  275.04 0.91 280.24 2.53 ;
      RECT  282.18 0.91 286.19 2.53 ;
      RECT  288.13 0.91 296.9 2.53 ;
      RECT  298.84 0.91 299.28 2.53 ;
      RECT  315.5 0.91 326.65 2.53 ;
      RECT  329.78 0.91 344.5 2.53 ;
      RECT  346.44 0.91 359.97 2.53 ;
      RECT  361.91 0.91 373.06 2.53 ;
      RECT  7.73 2.53 12.05 7.73 ;
      RECT  7.73 352.39 12.05 356.83 ;
      RECT  12.05 2.53 127.92 7.73 ;
      RECT  12.05 7.73 127.92 352.39 ;
      RECT  12.05 352.39 127.92 356.83 ;
      RECT  129.86 2.53 413.52 7.73 ;
      RECT  129.86 7.73 413.52 352.39 ;
      RECT  129.86 352.39 413.52 356.83 ;
      RECT  413.52 2.53 417.84 7.73 ;
      RECT  413.52 352.39 417.84 356.83 ;
      RECT  0.91 0.91 1.78 1.78 ;
      RECT  0.91 1.78 1.78 2.53 ;
      RECT  1.78 0.91 6.1 1.78 ;
      RECT  6.1 0.91 47.0 1.78 ;
      RECT  6.1 1.78 47.0 2.53 ;
      RECT  0.91 2.53 1.78 7.73 ;
      RECT  6.1 2.53 7.73 7.73 ;
      RECT  0.91 7.73 1.78 352.39 ;
      RECT  6.1 7.73 7.73 352.39 ;
      RECT  0.91 352.39 1.78 356.83 ;
      RECT  6.1 352.39 7.73 356.83 ;
      RECT  375.0 0.91 419.47 1.78 ;
      RECT  375.0 1.78 419.47 2.53 ;
      RECT  419.47 0.91 423.79 1.78 ;
      RECT  423.79 0.91 424.66 1.78 ;
      RECT  423.79 1.78 424.66 2.53 ;
      RECT  417.84 2.53 419.47 7.73 ;
      RECT  423.79 2.53 424.66 7.73 ;
      RECT  417.84 7.73 419.47 352.39 ;
      RECT  423.79 7.73 424.66 352.39 ;
      RECT  417.84 352.39 419.47 356.83 ;
      RECT  423.79 352.39 424.66 356.83 ;
   END
END    conv2_wm_sram_16_200_sky130A
END    LIBRARY
