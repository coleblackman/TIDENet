VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO conv2_rm_sram_16_288_sky130A
   CLASS BLOCK ;
   SIZE 432.71 BY 474.36 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  129.71 0.0 130.45 1.93 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  142.8 0.0 143.54 1.93 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  157.08 0.0 157.82 1.93 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  170.17 0.0 170.91 1.93 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  183.26 0.0 184.0 1.93 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  195.16 0.0 195.9 1.93 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  209.44 0.0 210.18 1.93 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  222.53 0.0 223.27 1.93 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  235.62 0.0 236.36 1.93 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  248.71 0.0 249.45 1.93 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  261.8 0.0 262.54 1.93 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  274.89 0.0 275.63 1.93 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  287.98 0.0 288.72 1.93 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  301.07 0.0 301.81 1.93 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  314.16 0.0 314.9 1.93 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  328.44 0.0 329.18 1.93 ;
      END
   END din0[15]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  103.53 0.0 104.27 1.93 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  116.62 0.0 117.36 1.93 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 183.26 1.93 184.0 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 184.45 1.93 185.19 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 190.4 1.93 191.14 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 192.78 1.93 193.52 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 199.92 1.93 200.66 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 201.11 1.93 201.85 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 207.06 1.93 207.8 ;
      END
   END addr0[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 29.75 1.93 30.49 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.0 33.32 1.93 34.06 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  48.79 0.0 49.53 1.93 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  159.46 0.0 160.2 1.93 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  176.12 0.0 176.86 1.93 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  192.78 0.0 193.52 1.93 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  208.25 0.0 208.99 1.93 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  223.72 0.0 224.46 1.93 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  236.81 0.0 237.55 1.93 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  255.85 0.0 256.59 1.93 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  272.51 0.0 273.25 1.93 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  289.17 0.0 289.91 1.93 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  303.45 0.0 304.19 1.93 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  320.11 0.0 320.85 1.93 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  337.96 0.0 338.7 1.93 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  352.24 0.0 352.98 1.93 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  367.71 0.0 368.45 1.93 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  384.37 0.0 385.11 1.93 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  430.78 35.7 432.71 36.44 ;
      END
   END dout0[15]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m4 ;
         RECT  8.33 8.33 11.45 468.41 ;
         LAYER m3 ;
         RECT  8.33 465.29 424.38 468.41 ;
         LAYER m4 ;
         RECT  421.26 8.33 424.38 468.41 ;
         LAYER m3 ;
         RECT  8.33 8.33 424.38 11.45 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m4 ;
         RECT  2.38 2.38 5.5 474.36 ;
         LAYER m4 ;
         RECT  427.21 2.38 430.33 474.36 ;
         LAYER m3 ;
         RECT  2.38 471.24 430.33 474.36 ;
         LAYER m3 ;
         RECT  2.38 2.38 430.33 5.5 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  0.91 0.91 431.8 473.45 ;
   LAYER  m2 ;
      RECT  0.91 0.91 431.8 473.45 ;
   LAYER  m3 ;
      RECT  2.83 182.36 431.8 184.9 ;
      RECT  0.91 186.09 2.83 189.5 ;
      RECT  0.91 194.42 2.83 199.02 ;
      RECT  0.91 202.75 2.83 206.16 ;
      RECT  0.91 31.39 2.83 32.42 ;
      RECT  0.91 34.96 2.83 182.36 ;
      RECT  2.83 34.8 429.88 37.34 ;
      RECT  2.83 37.34 429.88 182.36 ;
      RECT  429.88 37.34 431.8 182.36 ;
      RECT  2.83 184.9 7.43 464.39 ;
      RECT  2.83 464.39 7.43 469.31 ;
      RECT  7.43 184.9 425.28 464.39 ;
      RECT  425.28 184.9 431.8 464.39 ;
      RECT  425.28 464.39 431.8 469.31 ;
      RECT  2.83 7.43 7.43 12.35 ;
      RECT  2.83 12.35 7.43 34.8 ;
      RECT  7.43 12.35 425.28 34.8 ;
      RECT  425.28 7.43 429.88 12.35 ;
      RECT  425.28 12.35 429.88 34.8 ;
      RECT  0.91 208.7 1.48 470.34 ;
      RECT  0.91 470.34 1.48 473.45 ;
      RECT  1.48 208.7 2.83 470.34 ;
      RECT  2.83 469.31 7.43 470.34 ;
      RECT  7.43 469.31 425.28 470.34 ;
      RECT  425.28 469.31 431.23 470.34 ;
      RECT  431.23 469.31 431.8 470.34 ;
      RECT  431.23 470.34 431.8 473.45 ;
      RECT  0.91 0.91 1.48 1.48 ;
      RECT  0.91 1.48 1.48 6.4 ;
      RECT  0.91 6.4 1.48 28.85 ;
      RECT  1.48 0.91 2.83 1.48 ;
      RECT  1.48 6.4 2.83 28.85 ;
      RECT  429.88 0.91 431.23 1.48 ;
      RECT  429.88 6.4 431.23 34.8 ;
      RECT  431.23 0.91 431.8 1.48 ;
      RECT  431.23 1.48 431.8 6.4 ;
      RECT  431.23 6.4 431.8 34.8 ;
      RECT  2.83 0.91 7.43 1.48 ;
      RECT  2.83 6.4 7.43 7.43 ;
      RECT  7.43 0.91 425.28 1.48 ;
      RECT  7.43 6.4 425.28 7.43 ;
      RECT  425.28 0.91 429.88 1.48 ;
      RECT  425.28 6.4 429.88 7.43 ;
   LAYER  m4 ;
      RECT  129.11 2.53 131.05 473.45 ;
      RECT  131.05 0.91 142.2 2.53 ;
      RECT  144.14 0.91 156.48 2.53 ;
      RECT  210.78 0.91 221.93 2.53 ;
      RECT  276.23 0.91 287.38 2.53 ;
      RECT  104.87 0.91 116.02 2.53 ;
      RECT  117.96 0.91 129.11 2.53 ;
      RECT  50.13 0.91 102.93 2.53 ;
      RECT  158.42 0.91 158.86 2.53 ;
      RECT  160.8 0.91 169.57 2.53 ;
      RECT  171.51 0.91 175.52 2.53 ;
      RECT  177.46 0.91 182.66 2.53 ;
      RECT  184.6 0.91 192.18 2.53 ;
      RECT  194.12 0.91 194.56 2.53 ;
      RECT  196.5 0.91 207.65 2.53 ;
      RECT  225.06 0.91 235.02 2.53 ;
      RECT  238.15 0.91 248.11 2.53 ;
      RECT  250.05 0.91 255.25 2.53 ;
      RECT  257.19 0.91 261.2 2.53 ;
      RECT  263.14 0.91 271.91 2.53 ;
      RECT  273.85 0.91 274.29 2.53 ;
      RECT  290.51 0.91 300.47 2.53 ;
      RECT  302.41 0.91 302.85 2.53 ;
      RECT  304.79 0.91 313.56 2.53 ;
      RECT  315.5 0.91 319.51 2.53 ;
      RECT  321.45 0.91 327.84 2.53 ;
      RECT  329.78 0.91 337.36 2.53 ;
      RECT  339.3 0.91 351.64 2.53 ;
      RECT  353.58 0.91 367.11 2.53 ;
      RECT  369.05 0.91 383.77 2.53 ;
      RECT  7.73 2.53 12.05 7.73 ;
      RECT  7.73 469.01 12.05 473.45 ;
      RECT  12.05 2.53 129.11 7.73 ;
      RECT  12.05 7.73 129.11 469.01 ;
      RECT  12.05 469.01 129.11 473.45 ;
      RECT  131.05 2.53 420.66 7.73 ;
      RECT  131.05 7.73 420.66 469.01 ;
      RECT  131.05 469.01 420.66 473.45 ;
      RECT  420.66 2.53 424.98 7.73 ;
      RECT  420.66 469.01 424.98 473.45 ;
      RECT  0.91 0.91 1.78 1.78 ;
      RECT  0.91 1.78 1.78 2.53 ;
      RECT  1.78 0.91 6.1 1.78 ;
      RECT  6.1 0.91 48.19 1.78 ;
      RECT  6.1 1.78 48.19 2.53 ;
      RECT  0.91 2.53 1.78 7.73 ;
      RECT  6.1 2.53 7.73 7.73 ;
      RECT  0.91 7.73 1.78 469.01 ;
      RECT  6.1 7.73 7.73 469.01 ;
      RECT  0.91 469.01 1.78 473.45 ;
      RECT  6.1 469.01 7.73 473.45 ;
      RECT  385.71 0.91 426.61 1.78 ;
      RECT  385.71 1.78 426.61 2.53 ;
      RECT  426.61 0.91 430.93 1.78 ;
      RECT  430.93 0.91 431.8 1.78 ;
      RECT  430.93 1.78 431.8 2.53 ;
      RECT  424.98 2.53 426.61 7.73 ;
      RECT  430.93 2.53 431.8 7.73 ;
      RECT  424.98 7.73 426.61 469.01 ;
      RECT  430.93 7.73 431.8 469.01 ;
      RECT  424.98 469.01 426.61 473.45 ;
      RECT  430.93 469.01 431.8 473.45 ;
   END
END    conv2_rm_sram_16_288_sky130A
END    LIBRARY
